magic
tech scmos
timestamp 1383052641
<< metal1 >>
rect 1553 696 1563 699
rect 1546 687 1563 690
rect 2328 581 2335 584
rect 2328 468 2335 471
rect 2339 468 2362 471
rect 2339 458 2356 461
rect 575 349 578 382
rect 582 355 585 416
rect 2328 355 2335 358
rect 582 352 1187 355
rect 2339 355 2375 358
rect 575 346 1181 349
rect 1178 271 1181 346
rect 1184 278 1187 352
rect 2339 345 2369 348
rect 2328 282 2409 285
rect 1184 275 2376 278
rect 1178 268 2369 271
rect 1174 261 2363 264
rect 1166 254 2356 257
<< m2contact >>
rect 1563 696 1567 700
rect 1563 687 1567 691
rect 2335 580 2339 584
rect 2335 467 2339 471
rect 2362 467 2366 471
rect 2356 457 2360 461
rect 581 416 585 420
rect 575 382 579 386
rect 2335 354 2339 358
rect 2375 354 2379 358
rect 2369 344 2373 348
rect 2324 281 2328 285
rect 2376 274 2380 278
rect 2369 267 2373 271
rect 1170 261 1174 265
rect 2363 260 2367 264
rect 1162 254 1166 258
rect 2356 253 2360 257
<< metal2 >>
rect 1567 696 2393 699
rect 1567 687 2387 690
rect 2339 581 2353 584
rect 2339 571 2347 574
rect 578 416 581 420
rect 1165 303 1173 307
rect 1162 258 1165 276
rect 1170 265 1173 303
rect 1758 288 2327 291
rect 2324 285 2327 288
rect 2344 229 2347 571
rect 2334 225 2347 229
rect 2350 194 2353 581
rect 2357 257 2360 457
rect 2363 264 2366 467
rect 2370 271 2373 344
rect 2376 278 2379 354
rect 2338 190 2353 194
rect 2276 81 2277 82
rect 2384 81 2387 687
rect 2276 77 2387 81
rect 2390 16 2393 696
rect 1570 13 2393 16
use tree  tree_1
timestamp 1383046086
transform -1 0 2340 0 -1 620
box -2 -116 2352 334
use tree  tree_0
timestamp 1383046086
transform 1 0 -13 0 1 110
box -2 -116 2352 334
<< end >>
