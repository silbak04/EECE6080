magic
tech scmos
timestamp 1384231894
<< nwell >>
rect 20 739 280 999
rect 17 428 283 652
rect -3 247 303 329
rect -3 10 11 247
rect 289 10 303 247
rect -3 -4 303 10
<< pwell >>
rect -3 655 303 672
rect -3 425 14 655
rect 286 425 303 655
rect -3 339 303 425
rect 11 10 289 247
<< ntransistor >>
rect 38 215 138 218
rect 162 215 262 218
rect 38 170 138 173
rect 38 149 138 152
rect 162 170 262 173
rect 162 149 262 152
rect 38 105 138 108
rect 38 84 138 87
rect 162 105 262 108
rect 162 84 262 87
rect 38 40 138 43
rect 162 40 262 43
<< ndiffusion >>
rect 38 226 138 227
rect 38 222 41 226
rect 95 222 138 226
rect 38 218 138 222
rect 162 226 262 227
rect 162 222 205 226
rect 259 222 262 226
rect 162 218 262 222
rect 38 199 138 215
rect 38 195 56 199
rect 120 195 138 199
rect 38 193 138 195
rect 38 189 56 193
rect 120 189 138 193
rect 38 173 138 189
rect 38 166 138 170
rect 38 162 41 166
rect 120 162 138 166
rect 38 160 138 162
rect 38 156 41 160
rect 120 156 138 160
rect 38 152 138 156
rect 38 133 138 149
rect 38 124 56 133
rect 120 124 138 133
rect 38 108 138 124
rect 162 199 262 215
rect 162 195 180 199
rect 244 195 262 199
rect 162 193 262 195
rect 162 189 180 193
rect 244 189 262 193
rect 162 173 262 189
rect 162 166 262 170
rect 162 162 180 166
rect 259 162 262 166
rect 162 160 262 162
rect 162 156 180 160
rect 259 156 262 160
rect 162 152 262 156
rect 38 101 138 105
rect 38 97 41 101
rect 120 97 138 101
rect 38 95 138 97
rect 38 91 41 95
rect 120 91 138 95
rect 38 87 138 91
rect 38 68 138 84
rect 38 59 56 68
rect 120 59 138 68
rect 38 43 138 59
rect 162 133 262 149
rect 162 124 180 133
rect 244 124 262 133
rect 162 108 262 124
rect 162 101 262 105
rect 162 97 180 101
rect 259 97 262 101
rect 162 95 262 97
rect 162 91 180 95
rect 259 91 262 95
rect 162 87 262 91
rect 162 68 262 84
rect 162 59 180 68
rect 244 59 262 68
rect 162 43 262 59
rect 38 36 138 40
rect 38 32 41 36
rect 95 32 138 36
rect 38 31 138 32
rect 162 36 262 40
rect 162 32 205 36
rect 259 32 262 36
rect 162 31 262 32
<< ndcontact >>
rect 41 222 95 226
rect 205 222 259 226
rect 56 195 120 199
rect 56 189 120 193
rect 41 162 120 166
rect 41 156 120 160
rect 56 124 120 133
rect 180 195 244 199
rect 180 189 244 193
rect 180 162 259 166
rect 180 156 259 160
rect 41 97 120 101
rect 41 91 120 95
rect 56 59 120 68
rect 180 124 244 133
rect 180 97 259 101
rect 180 91 259 95
rect 180 59 244 68
rect 41 32 95 36
rect 205 32 259 36
<< psubstratepdiff >>
rect 0 668 300 669
rect 0 659 1 668
rect 95 659 204 668
rect 298 659 300 668
rect 0 658 300 659
rect 0 657 11 658
rect 0 423 1 657
rect 10 423 11 657
rect 289 657 300 658
rect 0 422 11 423
rect 289 423 290 657
rect 299 423 300 657
rect 289 422 300 423
rect 0 417 300 422
rect 0 413 143 417
rect 157 413 204 417
rect 298 413 300 417
rect 0 412 300 413
rect 0 408 2 412
rect 96 408 300 412
rect 0 407 300 408
rect 0 403 143 407
rect 157 403 204 407
rect 298 403 300 407
rect 0 402 300 403
rect 0 398 2 402
rect 96 398 300 402
rect 0 397 300 398
rect 0 393 143 397
rect 157 393 204 397
rect 298 393 300 397
rect 0 392 300 393
rect 0 388 2 392
rect 96 388 300 392
rect 0 387 300 388
rect 0 383 143 387
rect 157 383 204 387
rect 298 383 300 387
rect 0 382 300 383
rect 0 378 2 382
rect 96 378 300 382
rect 0 377 300 378
rect 0 373 143 377
rect 157 373 204 377
rect 298 373 300 377
rect 0 372 300 373
rect 0 368 2 372
rect 96 368 300 372
rect 0 367 300 368
rect 0 363 143 367
rect 157 363 204 367
rect 298 363 300 367
rect 0 362 300 363
rect 0 358 2 362
rect 96 358 300 362
rect 0 357 300 358
rect 0 353 143 357
rect 157 353 204 357
rect 298 353 300 357
rect 0 347 300 353
rect 0 343 2 347
rect 96 343 143 347
rect 157 343 204 347
rect 298 343 300 347
rect 0 342 300 343
rect 14 243 286 244
rect 14 240 202 243
rect 14 236 19 240
rect 98 236 202 240
rect 14 234 202 236
rect 281 234 286 243
rect 14 232 286 234
rect 14 28 24 232
rect 28 229 39 232
rect 28 29 30 229
rect 38 228 39 229
rect 98 229 202 232
rect 98 228 138 229
rect 38 227 138 228
rect 142 222 158 229
rect 142 218 145 222
rect 154 218 158 222
rect 162 228 202 229
rect 261 229 277 232
rect 261 228 262 229
rect 162 227 262 228
rect 142 214 158 218
rect 142 210 145 214
rect 154 210 158 214
rect 142 206 158 210
rect 142 202 145 206
rect 154 202 158 206
rect 142 134 158 202
rect 142 130 145 134
rect 154 130 158 134
rect 142 126 158 130
rect 142 122 145 126
rect 154 122 158 126
rect 142 62 158 122
rect 142 58 145 62
rect 154 58 158 62
rect 142 54 158 58
rect 142 50 145 54
rect 154 50 158 54
rect 142 46 158 50
rect 142 42 145 46
rect 154 42 158 46
rect 38 29 138 31
rect 142 38 158 42
rect 142 34 145 38
rect 154 34 158 38
rect 142 29 158 34
rect 162 29 262 31
rect 270 29 277 229
rect 28 28 277 29
rect 281 28 286 232
rect 14 26 286 28
rect 14 22 19 26
rect 98 22 202 26
rect 281 22 286 26
rect 14 13 286 22
<< nsubstratendiff >>
rect 20 648 280 649
rect 20 644 23 648
rect 277 644 280 648
rect 20 638 280 644
rect 20 634 23 638
rect 277 634 280 638
rect 20 628 280 634
rect 20 624 23 628
rect 277 624 280 628
rect 20 618 280 624
rect 20 614 23 618
rect 277 614 280 618
rect 20 608 280 614
rect 20 604 23 608
rect 277 604 280 608
rect 20 598 280 604
rect 20 594 23 598
rect 277 594 280 598
rect 20 588 280 594
rect 20 584 23 588
rect 277 584 280 588
rect 20 578 280 584
rect 20 574 23 578
rect 277 574 280 578
rect 20 568 280 574
rect 20 564 23 568
rect 277 564 280 568
rect 20 558 280 564
rect 20 554 23 558
rect 277 554 280 558
rect 20 548 280 554
rect 20 544 23 548
rect 277 544 280 548
rect 20 538 280 544
rect 20 534 23 538
rect 277 534 280 538
rect 20 528 280 534
rect 20 524 23 528
rect 277 524 280 528
rect 20 518 280 524
rect 20 514 23 518
rect 277 514 280 518
rect 20 508 280 514
rect 20 504 23 508
rect 277 504 280 508
rect 20 498 280 504
rect 20 494 23 498
rect 277 494 280 498
rect 20 488 280 494
rect 20 484 23 488
rect 277 484 280 488
rect 20 478 280 484
rect 20 474 23 478
rect 277 474 280 478
rect 20 468 280 474
rect 20 464 23 468
rect 277 464 280 468
rect 20 458 280 464
rect 20 454 23 458
rect 277 454 280 458
rect 20 448 280 454
rect 20 444 23 448
rect 277 444 280 448
rect 20 438 280 444
rect 20 434 23 438
rect 277 434 280 438
rect 20 431 280 434
rect 0 325 300 326
rect 0 321 3 325
rect 297 321 300 325
rect 0 315 300 321
rect 0 311 3 315
rect 297 311 300 315
rect 0 305 300 311
rect 0 301 3 305
rect 297 301 300 305
rect 0 295 300 301
rect 0 291 3 295
rect 297 291 300 295
rect 0 285 300 291
rect 0 281 3 285
rect 297 281 300 285
rect 0 275 300 281
rect 0 271 3 275
rect 297 271 300 275
rect 0 265 300 271
rect 0 261 3 265
rect 297 261 300 265
rect 0 255 300 261
rect 0 253 8 255
rect 0 4 2 253
rect 6 7 8 253
rect 292 253 300 255
rect 292 7 294 253
rect 6 6 294 7
rect 6 4 8 6
rect 0 2 8 4
rect 92 2 203 6
rect 292 4 294 6
rect 298 4 300 253
rect 292 2 300 4
rect 0 -1 300 2
<< psubstratepcontact >>
rect 1 659 95 668
rect 204 659 298 668
rect 1 423 10 657
rect 290 423 299 657
rect 143 413 157 417
rect 204 413 298 417
rect 2 408 96 412
rect 143 403 157 407
rect 204 403 298 407
rect 2 398 96 402
rect 143 393 157 397
rect 204 393 298 397
rect 2 388 96 392
rect 143 383 157 387
rect 204 383 298 387
rect 2 378 96 382
rect 143 373 157 377
rect 204 373 298 377
rect 2 368 96 372
rect 143 363 157 367
rect 204 363 298 367
rect 2 358 96 362
rect 143 353 157 357
rect 204 353 298 357
rect 2 343 96 347
rect 143 343 157 347
rect 204 343 298 347
rect 19 236 98 240
rect 202 234 281 243
rect 24 28 28 232
rect 39 228 98 232
rect 145 218 154 222
rect 202 228 261 232
rect 145 210 154 214
rect 145 202 154 206
rect 145 130 154 134
rect 145 122 154 126
rect 145 58 154 62
rect 145 50 154 54
rect 145 42 154 46
rect 145 34 154 38
rect 277 28 281 232
rect 19 22 98 26
rect 202 22 281 26
<< nsubstratencontact >>
rect 23 644 277 648
rect 23 634 277 638
rect 23 624 277 628
rect 23 614 277 618
rect 23 604 277 608
rect 23 594 277 598
rect 23 584 277 588
rect 23 574 277 578
rect 23 564 277 568
rect 23 554 277 558
rect 23 544 277 548
rect 23 534 277 538
rect 23 524 277 528
rect 23 514 277 518
rect 23 504 277 508
rect 23 494 277 498
rect 23 484 277 488
rect 23 474 277 478
rect 23 464 277 468
rect 23 454 277 458
rect 23 444 277 448
rect 23 434 277 438
rect 3 321 297 325
rect 3 311 297 315
rect 3 301 297 305
rect 3 291 297 295
rect 3 281 297 285
rect 3 271 297 275
rect 3 261 297 265
rect 2 4 6 253
rect 8 251 292 255
rect 8 2 92 6
rect 203 2 292 6
rect 294 4 298 253
<< polysilicon >>
rect 6 712 21 715
rect 24 712 39 715
rect 12 700 15 712
rect 24 709 27 712
rect 36 709 39 712
rect 24 706 39 709
rect 24 700 27 706
rect 36 700 39 706
rect 42 712 45 715
rect 42 709 51 712
rect 42 700 45 709
rect 48 706 51 709
rect 54 706 57 715
rect 48 703 57 706
rect 54 700 57 703
rect 60 712 63 715
rect 60 709 69 712
rect 60 700 63 709
rect 66 706 69 709
rect 72 706 75 715
rect 66 703 75 706
rect 72 700 75 703
rect 78 712 93 715
rect 96 712 111 715
rect 78 709 81 712
rect 96 709 99 712
rect 108 709 111 712
rect 78 706 93 709
rect 96 706 111 709
rect 190 706 205 709
rect 78 703 81 706
rect 78 700 93 703
rect 96 700 99 706
rect 105 700 108 706
rect 190 694 193 706
rect 196 700 199 706
rect 202 694 205 706
rect 208 706 223 709
rect 208 697 211 706
rect 220 697 223 706
rect 226 706 241 709
rect 244 706 259 709
rect 262 706 277 709
rect 226 703 229 706
rect 226 700 241 703
rect 238 697 241 700
rect 250 697 253 706
rect 262 703 265 706
rect 262 700 277 703
rect 274 697 277 700
rect 208 694 223 697
rect 226 694 241 697
rect 244 694 259 697
rect 262 694 277 697
rect 51 687 66 690
rect 69 687 84 690
rect 87 687 102 690
rect 51 678 54 687
rect 69 684 72 687
rect 87 684 90 687
rect 69 681 84 684
rect 87 681 102 684
rect 69 678 72 681
rect 99 678 102 681
rect 51 675 66 678
rect 69 675 84 678
rect 87 675 102 678
rect 31 216 38 218
rect 31 42 32 216
rect 36 215 38 216
rect 138 215 140 218
rect 36 173 37 215
rect 160 215 162 218
rect 262 216 269 218
rect 262 215 264 216
rect 36 170 38 173
rect 138 170 140 173
rect 36 152 37 170
rect 36 149 38 152
rect 138 149 140 152
rect 36 108 37 149
rect 263 173 264 215
rect 160 170 162 173
rect 262 170 264 173
rect 263 152 264 170
rect 160 149 162 152
rect 262 149 264 152
rect 36 105 38 108
rect 138 105 140 108
rect 36 87 37 105
rect 36 84 38 87
rect 138 84 140 87
rect 36 43 37 84
rect 263 108 264 149
rect 160 105 162 108
rect 262 105 264 108
rect 263 87 264 105
rect 160 84 162 87
rect 262 84 264 87
rect 36 42 38 43
rect 31 40 38 42
rect 138 40 140 43
rect 263 43 264 84
rect 160 40 162 43
rect 262 42 264 43
rect 268 42 269 216
rect 262 40 269 42
<< polycontact >>
rect 32 42 36 216
rect 264 42 268 216
<< metal1 >>
rect 20 996 280 999
rect 20 742 23 996
rect 277 742 280 996
rect 20 739 280 742
rect 62 729 238 739
rect 72 719 228 729
rect 82 709 218 719
rect 92 699 208 709
rect 0 668 99 669
rect 0 659 1 668
rect 95 659 99 668
rect 0 658 99 659
rect 0 657 10 658
rect 0 423 1 657
rect 102 649 198 699
rect 201 668 300 669
rect 201 659 204 668
rect 298 659 300 668
rect 201 658 300 659
rect 289 657 300 658
rect 50 648 280 649
rect 21 644 23 648
rect 277 644 280 648
rect 21 643 280 644
rect 21 639 23 643
rect 277 639 280 643
rect 21 638 280 639
rect 21 634 23 638
rect 277 634 280 638
rect 21 633 280 634
rect 21 629 23 633
rect 277 629 280 633
rect 21 628 280 629
rect 21 624 23 628
rect 277 624 280 628
rect 21 623 280 624
rect 21 619 23 623
rect 277 619 280 623
rect 21 618 280 619
rect 21 614 23 618
rect 277 614 280 618
rect 21 613 280 614
rect 21 609 23 613
rect 277 609 280 613
rect 21 608 280 609
rect 21 604 23 608
rect 277 604 280 608
rect 21 603 280 604
rect 21 599 23 603
rect 277 599 280 603
rect 21 598 280 599
rect 21 594 23 598
rect 277 594 280 598
rect 21 593 280 594
rect 21 589 23 593
rect 277 589 280 593
rect 21 588 280 589
rect 21 584 23 588
rect 277 584 280 588
rect 21 583 280 584
rect 21 579 23 583
rect 277 579 280 583
rect 21 578 280 579
rect 21 574 23 578
rect 277 574 280 578
rect 21 573 280 574
rect 21 569 23 573
rect 277 569 280 573
rect 21 568 280 569
rect 21 564 23 568
rect 277 564 280 568
rect 21 563 280 564
rect 21 559 23 563
rect 277 559 280 563
rect 21 558 280 559
rect 21 554 23 558
rect 277 554 280 558
rect 21 553 280 554
rect 21 549 23 553
rect 277 549 280 553
rect 21 548 280 549
rect 21 544 23 548
rect 277 544 280 548
rect 21 543 280 544
rect 21 539 23 543
rect 277 539 280 543
rect 21 538 280 539
rect 21 534 23 538
rect 277 534 280 538
rect 21 533 280 534
rect 21 529 23 533
rect 277 529 280 533
rect 21 528 280 529
rect 21 524 23 528
rect 277 524 280 528
rect 21 523 280 524
rect 21 519 23 523
rect 277 519 280 523
rect 21 518 280 519
rect 21 514 23 518
rect 277 514 280 518
rect 21 513 280 514
rect 21 509 23 513
rect 277 509 280 513
rect 21 508 280 509
rect 21 504 23 508
rect 277 504 280 508
rect 21 503 280 504
rect 21 499 23 503
rect 277 499 280 503
rect 21 498 280 499
rect 21 494 23 498
rect 277 494 280 498
rect 21 493 280 494
rect 21 489 23 493
rect 277 489 280 493
rect 21 488 280 489
rect 21 484 23 488
rect 277 484 280 488
rect 21 483 280 484
rect 21 479 23 483
rect 277 479 280 483
rect 21 478 280 479
rect 21 474 23 478
rect 277 474 280 478
rect 21 473 280 474
rect 21 469 23 473
rect 277 469 280 473
rect 21 468 280 469
rect 21 464 23 468
rect 277 464 280 468
rect 21 463 280 464
rect 21 459 23 463
rect 277 459 280 463
rect 21 458 280 459
rect 21 454 23 458
rect 277 454 280 458
rect 21 453 280 454
rect 21 449 23 453
rect 277 449 280 453
rect 21 448 280 449
rect 21 444 23 448
rect 277 444 280 448
rect 21 443 280 444
rect 21 439 23 443
rect 277 439 280 443
rect 21 438 280 439
rect 21 434 23 438
rect 277 434 280 438
rect 21 432 280 434
rect 0 418 10 423
rect 102 423 198 432
rect 0 417 99 418
rect 0 413 2 417
rect 96 413 99 417
rect 0 412 99 413
rect 0 408 2 412
rect 96 408 99 412
rect 0 407 99 408
rect 0 403 2 407
rect 96 403 99 407
rect 0 402 99 403
rect 0 398 2 402
rect 96 398 99 402
rect 0 397 99 398
rect 0 393 2 397
rect 96 393 99 397
rect 0 392 99 393
rect 0 388 2 392
rect 96 388 99 392
rect 0 387 99 388
rect 0 383 2 387
rect 96 383 99 387
rect 0 382 99 383
rect 0 378 2 382
rect 96 378 99 382
rect 0 377 99 378
rect 0 373 2 377
rect 96 373 99 377
rect 0 372 99 373
rect 0 368 2 372
rect 96 368 99 372
rect 0 367 99 368
rect 0 363 2 367
rect 96 363 99 367
rect 0 362 99 363
rect 0 358 2 362
rect 96 358 99 362
rect 0 357 99 358
rect 0 348 2 357
rect 96 348 99 357
rect 0 347 99 348
rect 0 343 2 347
rect 96 343 99 347
rect 102 339 140 423
rect 143 417 157 420
rect 143 412 157 413
rect 143 407 157 408
rect 143 402 157 403
rect 143 397 157 398
rect 143 392 157 393
rect 143 387 157 388
rect 143 382 157 383
rect 143 377 157 378
rect 143 372 157 373
rect 143 367 157 368
rect 143 362 157 363
rect 143 357 157 358
rect 143 352 157 353
rect 143 347 157 348
rect 160 339 198 423
rect 289 423 290 657
rect 299 423 300 657
rect 289 418 300 423
rect 201 417 300 418
rect 201 413 204 417
rect 298 413 300 417
rect 201 412 300 413
rect 201 408 204 412
rect 298 408 300 412
rect 201 407 300 408
rect 201 403 204 407
rect 298 403 300 407
rect 201 402 300 403
rect 201 398 204 402
rect 298 398 300 402
rect 201 397 300 398
rect 201 393 204 397
rect 298 393 300 397
rect 201 392 300 393
rect 201 388 204 392
rect 298 388 300 392
rect 201 387 300 388
rect 201 383 204 387
rect 298 383 300 387
rect 201 382 300 383
rect 201 378 204 382
rect 298 378 300 382
rect 201 377 300 378
rect 201 373 204 377
rect 298 373 300 377
rect 201 372 300 373
rect 201 368 204 372
rect 298 368 300 372
rect 201 367 300 368
rect 201 363 204 367
rect 298 363 300 367
rect 201 362 300 363
rect 201 358 204 362
rect 298 358 300 362
rect 201 357 300 358
rect 201 353 204 357
rect 298 353 300 357
rect 201 352 300 353
rect 201 348 204 352
rect 298 348 300 352
rect 201 347 300 348
rect 201 343 204 347
rect 298 343 300 347
rect 102 325 198 339
rect 0 321 3 325
rect 297 321 300 325
rect 0 320 300 321
rect 0 316 3 320
rect 297 316 300 320
rect 0 315 300 316
rect 0 311 3 315
rect 297 311 300 315
rect 0 310 300 311
rect 0 306 3 310
rect 297 306 300 310
rect 0 305 300 306
rect 0 301 3 305
rect 297 301 300 305
rect 0 300 300 301
rect 0 296 3 300
rect 297 296 300 300
rect 0 295 300 296
rect 0 291 3 295
rect 297 291 300 295
rect 0 290 300 291
rect 0 286 3 290
rect 297 286 300 290
rect 0 285 300 286
rect 0 281 3 285
rect 297 281 300 285
rect 0 280 300 281
rect 0 276 3 280
rect 297 276 300 280
rect 0 275 300 276
rect 0 271 3 275
rect 297 271 300 275
rect 0 270 300 271
rect 0 266 3 270
rect 297 266 300 270
rect 0 265 300 266
rect 0 261 3 265
rect 297 261 300 265
rect 0 260 300 261
rect 0 256 8 260
rect 292 256 300 260
rect 0 255 300 256
rect 0 253 8 255
rect 0 4 2 253
rect 6 251 8 253
rect 292 253 300 255
rect 292 251 294 253
rect 6 250 294 251
rect 6 7 8 250
rect 14 240 99 245
rect 14 236 19 240
rect 98 236 99 240
rect 14 232 99 236
rect 14 227 24 232
rect 14 28 19 227
rect 23 28 24 227
rect 28 228 39 232
rect 98 228 99 232
rect 28 226 99 228
rect 28 222 41 226
rect 95 222 99 226
rect 28 216 99 222
rect 28 42 32 216
rect 36 214 99 216
rect 36 195 39 214
rect 53 210 57 214
rect 96 210 99 214
rect 102 229 198 250
rect 102 207 142 229
rect 36 193 53 195
rect 36 174 39 193
rect 56 199 142 207
rect 157 207 198 229
rect 201 243 286 245
rect 201 234 202 243
rect 281 234 286 243
rect 201 232 286 234
rect 201 228 202 232
rect 261 228 277 232
rect 201 227 277 228
rect 201 226 272 227
rect 201 222 205 226
rect 259 222 272 226
rect 201 216 272 222
rect 201 214 264 216
rect 201 210 204 214
rect 243 210 247 214
rect 157 199 244 207
rect 120 195 180 199
rect 56 193 244 195
rect 120 189 180 193
rect 56 181 244 189
rect 261 195 264 214
rect 247 193 264 195
rect 53 174 57 178
rect 116 174 120 178
rect 36 166 120 174
rect 36 162 41 166
rect 36 160 120 162
rect 36 156 41 160
rect 36 148 120 156
rect 36 109 39 148
rect 53 144 57 148
rect 116 144 120 148
rect 123 141 177 181
rect 180 174 184 178
rect 243 174 247 178
rect 261 174 264 193
rect 180 166 264 174
rect 259 162 264 166
rect 180 160 264 162
rect 259 156 264 160
rect 180 148 264 156
rect 180 144 184 148
rect 243 144 247 148
rect 56 137 244 141
rect 56 133 142 137
rect 120 124 142 133
rect 56 119 142 124
rect 157 133 244 137
rect 157 124 180 133
rect 157 119 244 124
rect 56 116 244 119
rect 53 109 57 113
rect 116 109 120 113
rect 36 101 120 109
rect 36 97 41 101
rect 36 95 120 97
rect 36 91 41 95
rect 36 83 120 91
rect 36 44 39 83
rect 53 79 57 83
rect 116 79 120 83
rect 123 76 177 116
rect 180 109 184 113
rect 243 109 247 113
rect 261 109 264 148
rect 180 101 264 109
rect 259 97 264 101
rect 180 95 264 97
rect 259 91 264 95
rect 180 83 264 91
rect 180 79 184 83
rect 243 79 247 83
rect 56 69 244 76
rect 56 68 142 69
rect 120 59 142 68
rect 157 68 244 69
rect 56 51 142 59
rect 53 44 57 48
rect 96 44 99 48
rect 36 42 99 44
rect 28 36 99 42
rect 28 32 41 36
rect 95 32 99 36
rect 28 28 39 32
rect 98 28 99 32
rect 14 26 99 28
rect 14 22 19 26
rect 98 22 99 26
rect 14 21 99 22
rect 14 17 19 21
rect 98 17 99 21
rect 14 13 99 17
rect 102 27 142 51
rect 157 59 180 68
rect 157 51 244 59
rect 157 27 198 51
rect 6 6 99 7
rect 6 4 8 6
rect 0 2 8 4
rect 92 2 99 6
rect 0 -1 99 2
rect 102 -1 198 27
rect 201 44 204 48
rect 243 44 247 48
rect 261 44 264 83
rect 201 42 264 44
rect 268 42 272 216
rect 201 36 272 42
rect 201 32 205 36
rect 259 32 272 36
rect 201 28 202 32
rect 261 28 272 32
rect 276 28 277 227
rect 281 28 286 232
rect 201 26 286 28
rect 201 22 202 26
rect 281 22 286 26
rect 201 21 286 22
rect 201 17 202 21
rect 281 17 286 21
rect 201 13 286 17
rect 292 7 294 250
rect 201 6 294 7
rect 201 2 203 6
rect 292 4 294 6
rect 298 4 300 253
rect 292 2 300 4
rect 201 -1 300 2
<< m2contact >>
rect 23 639 277 643
rect 23 629 277 633
rect 23 619 277 623
rect 23 609 277 613
rect 23 599 277 603
rect 23 589 277 593
rect 23 579 277 583
rect 23 569 277 573
rect 23 559 277 563
rect 23 549 277 553
rect 23 539 277 543
rect 23 529 277 533
rect 23 519 277 523
rect 23 509 277 513
rect 23 499 277 503
rect 23 489 277 493
rect 23 479 277 483
rect 23 469 277 473
rect 23 459 277 463
rect 23 449 277 453
rect 23 439 277 443
rect 2 413 96 417
rect 2 403 96 407
rect 2 393 96 397
rect 2 383 96 387
rect 2 373 96 377
rect 2 363 96 367
rect 2 348 96 357
rect 143 408 157 412
rect 143 398 157 402
rect 143 388 157 392
rect 143 378 157 382
rect 143 368 157 372
rect 143 358 157 362
rect 143 348 157 352
rect 204 408 298 412
rect 204 398 298 402
rect 204 388 298 392
rect 204 378 298 382
rect 204 368 298 372
rect 204 358 298 362
rect 204 348 298 352
rect 3 316 297 320
rect 3 306 297 310
rect 3 296 297 300
rect 3 286 297 290
rect 3 276 297 280
rect 3 266 297 270
rect 8 256 292 260
rect 19 28 23 227
rect 39 195 53 214
rect 57 210 96 214
rect 39 174 53 193
rect 145 222 154 226
rect 145 214 154 218
rect 145 206 154 210
rect 204 210 243 214
rect 247 195 261 214
rect 57 174 116 178
rect 39 109 53 148
rect 57 144 116 148
rect 184 174 243 178
rect 247 174 261 193
rect 184 144 243 148
rect 145 126 154 130
rect 57 109 116 113
rect 39 44 53 83
rect 57 79 116 83
rect 184 109 243 113
rect 247 109 261 148
rect 184 79 243 83
rect 57 44 96 48
rect 39 28 98 32
rect 19 17 98 21
rect 145 62 154 66
rect 145 54 154 58
rect 145 46 154 50
rect 145 38 154 42
rect 145 30 154 34
rect 204 44 243 48
rect 247 44 261 83
rect 202 28 261 32
rect 272 28 276 227
rect 202 17 281 21
<< metal2 >>
rect 20 996 280 999
rect 20 742 23 996
rect 277 742 280 996
rect 20 739 280 742
rect 0 643 300 669
rect 0 639 23 643
rect 277 639 300 643
rect 0 633 300 639
rect 0 629 23 633
rect 277 629 300 633
rect 0 623 300 629
rect 0 619 23 623
rect 277 619 300 623
rect 0 613 300 619
rect 0 609 23 613
rect 277 609 300 613
rect 0 603 300 609
rect 0 599 23 603
rect 277 599 300 603
rect 0 593 300 599
rect 0 589 23 593
rect 277 589 300 593
rect 0 583 300 589
rect 0 579 23 583
rect 277 579 300 583
rect 0 573 300 579
rect 0 569 23 573
rect 277 569 300 573
rect 0 563 300 569
rect 0 559 23 563
rect 277 559 300 563
rect 0 553 300 559
rect 0 549 23 553
rect 277 549 300 553
rect 0 543 300 549
rect 0 539 23 543
rect 277 539 300 543
rect 0 533 300 539
rect 0 529 23 533
rect 277 529 300 533
rect 0 523 300 529
rect 0 519 23 523
rect 277 519 300 523
rect 0 513 300 519
rect 0 509 23 513
rect 277 509 300 513
rect 0 503 300 509
rect 0 499 23 503
rect 277 499 300 503
rect 0 493 300 499
rect 0 489 23 493
rect 277 489 300 493
rect 0 483 300 489
rect 0 479 23 483
rect 277 479 300 483
rect 0 473 300 479
rect 0 469 23 473
rect 277 469 300 473
rect 0 463 300 469
rect 0 459 23 463
rect 277 459 300 463
rect 0 453 300 459
rect 0 449 23 453
rect 277 449 300 453
rect 0 443 300 449
rect 0 439 23 443
rect 277 439 300 443
rect 0 417 300 423
rect 0 413 2 417
rect 96 413 300 417
rect 0 412 300 413
rect 0 408 143 412
rect 157 408 204 412
rect 298 408 300 412
rect 0 407 300 408
rect 0 403 2 407
rect 96 403 300 407
rect 0 402 300 403
rect 0 398 143 402
rect 157 398 204 402
rect 298 398 300 402
rect 0 397 300 398
rect 0 393 2 397
rect 96 393 300 397
rect 0 392 300 393
rect 0 388 143 392
rect 157 388 204 392
rect 298 388 300 392
rect 0 387 300 388
rect 0 383 2 387
rect 96 383 300 387
rect 0 382 300 383
rect 0 378 143 382
rect 157 378 204 382
rect 298 378 300 382
rect 0 377 300 378
rect 0 373 2 377
rect 96 373 300 377
rect 0 372 300 373
rect 0 368 143 372
rect 157 368 204 372
rect 298 368 300 372
rect 0 367 300 368
rect 0 363 2 367
rect 96 363 300 367
rect 0 362 300 363
rect 0 358 143 362
rect 157 358 204 362
rect 298 358 300 362
rect 0 357 300 358
rect 0 348 2 357
rect 96 352 300 357
rect 96 348 143 352
rect 157 348 204 352
rect 298 348 300 352
rect 0 343 300 348
rect 0 320 300 325
rect 0 316 3 320
rect 297 316 300 320
rect 0 310 300 316
rect 0 306 3 310
rect 297 306 300 310
rect 0 300 300 306
rect 0 296 3 300
rect 297 296 300 300
rect 0 290 300 296
rect 0 286 3 290
rect 297 286 300 290
rect 0 280 300 286
rect 0 276 3 280
rect 297 276 300 280
rect 0 270 300 276
rect 0 266 3 270
rect 297 266 300 270
rect 0 260 300 266
rect 0 256 8 260
rect 292 256 300 260
rect 0 245 300 256
rect 0 227 300 229
rect 0 28 19 227
rect 23 226 272 227
rect 23 222 145 226
rect 154 222 272 226
rect 23 218 272 222
rect 23 214 145 218
rect 154 214 272 218
rect 23 195 39 214
rect 53 210 57 214
rect 96 210 204 214
rect 243 210 247 214
rect 53 206 145 210
rect 154 206 247 210
rect 53 195 247 206
rect 261 195 272 214
rect 23 193 272 195
rect 23 174 39 193
rect 53 178 247 193
rect 53 174 57 178
rect 116 174 184 178
rect 243 174 247 178
rect 261 174 272 193
rect 23 148 272 174
rect 23 109 39 148
rect 53 144 57 148
rect 116 144 184 148
rect 243 144 247 148
rect 53 130 247 144
rect 53 126 145 130
rect 154 126 247 130
rect 53 113 247 126
rect 53 109 57 113
rect 116 109 184 113
rect 243 109 247 113
rect 261 109 272 148
rect 23 83 272 109
rect 23 44 39 83
rect 53 79 57 83
rect 116 79 184 83
rect 243 79 247 83
rect 53 66 247 79
rect 53 62 145 66
rect 154 62 247 66
rect 53 58 247 62
rect 53 54 145 58
rect 154 54 247 58
rect 53 50 247 54
rect 53 48 145 50
rect 53 44 57 48
rect 96 46 145 48
rect 154 48 247 50
rect 154 46 204 48
rect 96 44 204 46
rect 243 44 247 48
rect 261 44 272 83
rect 23 42 272 44
rect 23 38 145 42
rect 154 38 272 42
rect 23 34 272 38
rect 23 32 145 34
rect 23 28 39 32
rect 98 30 145 32
rect 154 32 272 34
rect 154 30 202 32
rect 98 28 202 30
rect 261 28 272 32
rect 276 28 300 227
rect 0 21 300 28
rect 0 17 19 21
rect 98 17 202 21
rect 281 17 300 21
rect 0 6 300 17
rect 0 -1 98 6
rect 202 -1 300 6
<< pad >>
rect 23 742 277 996
<< labels >>
rlabel metal1 150 -1 150 -1 8 Vdd
rlabel metal2 140 126 140 126 6 gnd:2
<< end >>
