magic
tech scmos
timestamp 1382957000
<< metal1 >>
rect 37 36 51 40
rect 47 26 51 36
use MUX2X1  MUX2X1_0
timestamp 1053021328
transform 1 0 3 0 1 3
box -5 -3 53 105
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 45 0 1 3
box -9 -3 26 105
<< end >>
