magic
tech scmos
timestamp 1383894975
<< nwell >>
rect 920 2564 948 2570
<< metal1 >>
rect 72 2664 100 2670
rect 920 2664 948 2670
rect 1771 2664 1806 2670
rect -763 2560 -760 2648
rect 30 2621 46 2624
rect 83 2624 87 2652
rect 930 2624 934 2652
rect 76 2620 87 2624
rect 878 2621 892 2624
rect 924 2620 934 2624
rect 1726 2621 1741 2624
rect -763 2557 -756 2560
rect -759 1894 -756 2557
rect -753 2538 -748 2569
rect 70 2564 98 2570
rect 920 2564 948 2570
rect 151 2545 213 2549
rect -697 2541 -639 2545
rect -697 2533 -693 2541
rect -731 1894 -727 1916
rect -700 1900 -697 1917
rect -686 1904 -648 1907
rect -700 1897 -654 1900
rect -759 1891 -755 1894
rect -758 1887 -755 1891
rect -731 1890 -661 1894
rect -758 1884 -668 1887
rect -671 1831 -668 1884
rect -665 1840 -661 1890
rect -657 1849 -654 1897
rect -651 1855 -648 1904
rect -643 1862 -639 2541
rect 151 2534 155 2545
rect -451 1920 -447 1927
rect -643 1858 -628 1862
rect -651 1852 -621 1855
rect -657 1848 -640 1849
rect -657 1846 -643 1848
rect -665 1836 -646 1840
rect -624 1838 -621 1852
rect -671 1827 -614 1831
rect -618 1823 -614 1827
rect -608 1830 -604 1904
rect 31 1906 35 1928
rect 209 1913 213 2545
rect 933 2541 1003 2545
rect 1032 2541 1059 2544
rect 933 2519 937 2541
rect 999 2534 1003 2541
rect 933 2392 937 2414
rect 397 1920 401 1928
rect 882 1927 883 1929
rect 209 1909 210 1913
rect -578 1844 -575 1904
rect 31 1902 371 1906
rect -451 1892 -447 1901
rect -126 1893 240 1897
rect -126 1892 -122 1893
rect -451 1888 -122 1892
rect 269 1888 272 1894
rect 367 1893 371 1902
rect 367 1890 486 1893
rect 506 1894 535 1897
rect 879 1895 883 1927
rect 933 1913 937 1923
rect 911 1909 937 1913
rect 965 1908 969 1917
rect 1018 1908 1021 1918
rect 1028 1908 1031 1930
rect 1056 1901 1059 2541
rect 1249 1922 1253 1928
rect 1151 1903 1225 1904
rect 894 1899 1059 1901
rect 891 1898 1059 1899
rect 1063 1900 1225 1903
rect 1063 1895 1066 1900
rect 1221 1897 1225 1900
rect 879 1892 1066 1895
rect 367 1889 490 1890
rect 509 1889 876 1890
rect 1088 1889 1092 1893
rect -33 1884 272 1888
rect 509 1886 1092 1889
rect 509 1883 513 1886
rect 876 1885 1090 1886
rect -358 1876 118 1880
rect -404 1869 -323 1872
rect -316 1864 107 1868
rect -316 1862 -312 1864
rect -567 1858 -312 1862
rect -140 1857 107 1860
rect -140 1854 -137 1857
rect -567 1851 -137 1854
rect 71 1845 103 1848
rect -578 1841 -362 1844
rect -365 1838 -362 1841
rect -365 1835 105 1838
rect -608 1826 105 1830
rect -618 1820 -589 1823
rect -593 1816 -589 1820
rect -593 1771 -590 1786
rect 114 1776 118 1876
rect 121 1856 124 1877
rect 139 1868 143 1877
rect 132 1864 143 1868
rect 155 1867 158 1877
rect 420 1879 513 1883
rect 540 1882 873 1883
rect 1119 1882 1122 1893
rect 540 1880 1122 1882
rect 869 1879 1122 1880
rect 172 1868 175 1877
rect 214 1864 218 1877
rect 525 1871 927 1875
rect 525 1864 529 1871
rect 214 1860 529 1864
rect 539 1867 921 1868
rect 539 1865 918 1867
rect 539 1856 542 1865
rect 121 1853 542 1856
rect 826 1860 915 1862
rect 826 1859 1233 1860
rect 826 1857 830 1859
rect 912 1857 1233 1859
rect 104 1772 118 1776
rect 126 1601 129 1845
rect 151 1821 154 1834
rect 826 1830 829 1853
rect 839 1826 843 1852
rect 1021 1851 1222 1854
rect 1021 1848 1025 1851
rect 1249 1847 1253 1903
rect 884 1800 888 1843
rect 1037 1842 1253 1847
rect 1258 1843 1261 1898
rect 1509 1857 1708 1860
rect 1504 1851 1701 1854
rect 1037 1836 1040 1842
rect 1643 1840 1715 1843
rect 1727 1837 1731 1927
rect 1755 1856 1786 1859
rect 1755 1850 1786 1853
rect 891 1770 894 1836
rect 898 1832 1040 1836
rect 1570 1834 1731 1837
rect 200 1739 219 1743
rect 200 1654 204 1739
rect 684 1684 720 1687
rect 884 1667 887 1684
rect 899 1673 903 1832
rect 1570 1829 1573 1834
rect 910 1826 1573 1829
rect 877 1664 887 1667
rect 824 1620 842 1624
rect 126 1598 145 1601
rect 142 1429 145 1598
rect 838 1539 842 1620
rect 846 1576 849 1621
rect 846 1573 856 1576
rect 836 1535 842 1539
rect 846 1508 849 1566
rect 836 1505 849 1508
rect 200 1501 219 1505
rect 142 1426 177 1429
rect 144 1347 148 1410
rect 144 1344 155 1347
rect 130 1301 143 1304
rect 104 1290 108 1294
rect 128 1290 143 1294
rect 116 1164 143 1167
rect 119 1133 143 1137
rect 151 1118 155 1344
rect 174 1317 177 1426
rect 194 1409 197 1451
rect 200 1420 204 1501
rect 853 1494 856 1573
rect 826 1491 856 1494
rect 686 1446 717 1449
rect 200 1416 207 1420
rect 194 1406 205 1409
rect 202 1389 205 1406
rect 202 1385 207 1389
rect 824 1382 845 1386
rect 183 1328 251 1331
rect 177 1182 180 1280
rect 162 1133 176 1137
rect 127 1114 155 1118
rect 127 1111 131 1114
rect 127 1107 135 1111
rect 101 1070 125 1073
rect -525 1044 -503 1048
rect -525 971 -520 1044
rect 114 1041 125 1044
rect 115 1010 125 1014
rect 132 980 135 1107
rect 183 1073 186 1328
rect 190 1284 193 1319
rect 841 1301 845 1382
rect 197 1263 220 1267
rect 191 1150 194 1220
rect 197 1182 201 1263
rect 677 1208 701 1211
rect 197 1178 205 1182
rect 858 1178 861 1357
rect 191 1147 205 1150
rect 822 1144 849 1148
rect 845 1098 849 1144
rect 330 1088 358 1091
rect 877 1091 880 1664
rect 887 1633 901 1637
rect 888 1515 901 1519
rect 888 1401 892 1515
rect 899 1424 902 1501
rect 910 1401 913 1826
rect 1553 1762 1560 1766
rect 939 1516 946 1520
rect 896 1144 911 1148
rect 815 1088 880 1091
rect 143 1070 186 1073
rect 142 1041 207 1044
rect 166 1025 217 1029
rect 166 1014 170 1025
rect 144 1010 170 1014
rect -607 967 -520 971
rect 127 976 135 980
rect 127 956 131 976
rect 838 972 841 1069
rect 933 1034 946 1038
rect 134 969 691 972
rect 134 963 137 969
rect 838 969 926 972
rect 909 959 921 962
rect -118 952 131 956
rect 773 952 830 956
rect 910 952 925 956
rect -343 924 -124 927
rect -343 914 -340 924
rect -233 903 -230 917
rect -224 905 -220 917
rect -127 907 -124 924
rect -118 921 -114 952
rect -97 943 156 947
rect 827 943 830 952
rect 845 943 920 948
rect -752 882 -746 898
rect -652 882 -646 893
rect -97 891 -94 943
rect 30 936 145 939
rect 12 915 15 936
rect 26 914 29 936
rect 152 930 156 943
rect 716 939 817 942
rect 163 936 719 939
rect 845 933 848 943
rect 751 930 848 933
rect 56 923 121 927
rect 152 926 261 930
rect 56 914 60 923
rect 117 921 121 923
rect 257 921 261 926
rect 274 924 601 928
rect 117 917 197 921
rect 257 917 625 921
rect 509 910 613 913
rect -67 903 135 907
rect -67 893 -63 903
rect -37 895 135 898
rect -224 879 -220 885
rect -222 878 -220 879
rect -769 336 -747 342
rect -769 142 -763 336
rect -37 258 -34 895
rect 88 887 132 890
rect 88 886 133 887
rect 88 857 92 886
rect 142 878 145 910
rect 169 900 172 910
rect 190 899 194 910
rect 622 904 625 917
rect 605 886 628 890
rect 751 887 754 930
rect 817 905 820 921
rect 827 905 830 921
rect 838 905 842 923
rect 874 912 877 932
rect 880 912 884 932
rect 917 927 920 943
rect 838 901 902 905
rect 906 901 909 905
rect 924 898 928 932
rect 933 921 938 1034
rect 949 969 979 972
rect 976 966 1676 969
rect 948 960 1668 963
rect 947 953 1640 957
rect 956 949 957 950
rect 956 946 979 949
rect 959 945 979 946
rect 955 939 1004 942
rect 946 935 982 936
rect 946 932 978 935
rect 963 925 1444 928
rect 933 918 1095 921
rect 933 917 1383 918
rect 1030 914 1383 917
rect 993 910 994 914
rect 781 894 928 898
rect 785 893 786 894
rect 624 879 628 886
rect 88 390 92 407
rect 22 260 26 273
rect 817 263 820 887
rect 990 879 994 910
rect 1472 879 1476 886
rect 937 396 941 409
rect 817 260 842 263
rect 870 261 874 272
rect 1665 264 1668 960
rect 1673 939 1676 966
rect 1684 961 1725 964
rect 1722 948 1725 961
rect 1752 949 1756 960
rect 1665 261 1679 264
rect -37 256 3 258
rect 22 256 88 260
rect 870 257 937 261
rect 1772 257 1778 276
rect 1792 264 1796 956
rect -37 255 6 256
rect 1772 251 1822 257
rect 79 236 100 242
rect 923 236 952 242
rect 1772 236 1778 251
rect 89 182 101 186
rect 89 176 93 182
rect 129 181 147 185
rect 937 182 949 186
rect 937 176 941 182
rect 977 181 995 184
rect 1792 182 1795 244
rect 1776 179 1795 182
rect -769 136 -750 142
rect 79 136 100 142
rect 928 136 949 142
<< m2contact >>
rect -763 2648 -759 2652
rect 46 2621 50 2625
rect 87 2648 91 2652
rect 934 2648 938 2652
rect 892 2620 896 2624
rect 1741 2621 1745 2625
rect -701 2513 -697 2517
rect -676 1930 -672 1934
rect -731 1916 -727 1920
rect -700 1917 -696 1921
rect -690 1904 -686 1908
rect 147 2513 151 2517
rect -455 1944 -451 1948
rect 27 1944 31 1948
rect 172 1930 176 1934
rect -451 1916 -447 1920
rect -608 1904 -604 1908
rect -628 1858 -624 1862
rect -643 1844 -639 1848
rect -646 1836 -642 1840
rect -624 1834 -620 1838
rect -578 1904 -574 1908
rect 1028 2541 1032 2545
rect 933 2515 937 2519
rect 995 2513 999 2517
rect 933 2414 937 2418
rect 933 2388 937 2392
rect 393 1944 397 1948
rect 875 1944 879 1948
rect 1027 1930 1031 1934
rect 397 1916 401 1920
rect 210 1909 214 1913
rect -451 1901 -447 1905
rect 240 1893 244 1897
rect 269 1894 273 1898
rect 486 1890 490 1894
rect 502 1893 506 1897
rect 535 1893 539 1897
rect 933 1923 937 1927
rect 965 1917 969 1921
rect 1017 1918 1021 1922
rect 911 1905 915 1909
rect 965 1904 969 1908
rect 1018 1904 1022 1908
rect 1027 1904 1031 1908
rect 890 1899 894 1903
rect 1241 1944 1245 1948
rect 1723 1944 1727 1948
rect 1249 1918 1253 1922
rect 1088 1893 1092 1897
rect -37 1884 -33 1888
rect 1119 1893 1123 1897
rect -362 1876 -358 1880
rect -408 1869 -404 1873
rect -323 1869 -319 1873
rect 107 1864 111 1868
rect -571 1858 -567 1862
rect 107 1857 111 1861
rect -571 1851 -567 1855
rect 67 1845 71 1849
rect 103 1845 107 1849
rect 105 1835 109 1839
rect 105 1826 109 1830
rect -593 1786 -589 1790
rect 84 1782 88 1786
rect 121 1877 125 1881
rect 139 1877 143 1881
rect 154 1877 158 1881
rect 128 1864 132 1868
rect 172 1877 176 1881
rect 214 1877 218 1881
rect 416 1879 420 1883
rect 536 1879 540 1883
rect 1221 1892 1225 1897
rect 1249 1903 1253 1907
rect 155 1863 159 1867
rect 172 1864 176 1868
rect 927 1871 931 1875
rect 918 1863 922 1867
rect 1233 1857 1237 1861
rect 826 1853 830 1857
rect 125 1845 129 1849
rect 150 1834 154 1838
rect 839 1852 843 1856
rect 826 1826 830 1830
rect 1222 1850 1226 1854
rect 839 1822 843 1826
rect 884 1843 888 1847
rect 1021 1844 1025 1848
rect 151 1817 155 1821
rect 1258 1898 1262 1902
rect 1505 1857 1509 1861
rect 1708 1856 1712 1860
rect 1500 1850 1504 1854
rect 1701 1850 1705 1854
rect 884 1796 888 1800
rect 891 1836 895 1840
rect 1258 1838 1263 1843
rect 1639 1840 1643 1844
rect 1715 1840 1719 1844
rect 1751 1856 1755 1860
rect 1751 1849 1755 1853
rect 891 1766 895 1770
rect 236 1743 240 1747
rect 680 1684 684 1688
rect 720 1684 724 1688
rect 884 1684 888 1688
rect 903 1673 907 1677
rect 204 1654 208 1658
rect 803 1624 807 1628
rect 846 1621 850 1625
rect 832 1535 836 1539
rect 846 1566 850 1570
rect 236 1505 240 1509
rect 832 1505 836 1509
rect 193 1451 197 1455
rect 144 1410 148 1414
rect 126 1301 130 1305
rect 143 1301 147 1305
rect 108 1290 112 1294
rect 124 1290 128 1294
rect 143 1290 147 1294
rect 83 1286 87 1290
rect 112 1164 116 1168
rect 143 1164 147 1168
rect 115 1133 119 1137
rect 143 1133 147 1137
rect 682 1446 686 1450
rect 717 1446 721 1450
rect 207 1416 211 1420
rect 207 1385 211 1389
rect 803 1386 807 1390
rect 174 1313 178 1317
rect 176 1280 180 1284
rect 176 1178 180 1182
rect 158 1133 162 1137
rect 176 1133 180 1137
rect 97 1070 101 1074
rect 125 1070 129 1074
rect -486 1040 -482 1044
rect 110 1041 114 1045
rect 125 1041 129 1045
rect 111 1010 115 1014
rect 125 1010 129 1014
rect 139 1070 143 1074
rect 251 1327 255 1331
rect 189 1319 193 1323
rect 857 1357 861 1361
rect 841 1297 845 1301
rect 189 1280 193 1284
rect 236 1267 240 1271
rect 190 1220 194 1224
rect 819 1240 823 1244
rect 673 1208 677 1212
rect 701 1208 705 1212
rect 205 1178 209 1182
rect 858 1174 862 1178
rect 205 1147 209 1151
rect 801 1148 805 1152
rect 218 1119 222 1123
rect 845 1094 849 1098
rect 326 1088 330 1092
rect 358 1088 362 1092
rect 811 1088 815 1092
rect 883 1633 887 1637
rect 901 1633 905 1637
rect 901 1515 905 1519
rect 899 1501 903 1505
rect 899 1420 903 1424
rect 892 1401 896 1405
rect 1532 1766 1536 1770
rect 1560 1762 1564 1766
rect 943 1752 947 1756
rect 963 1520 967 1524
rect 916 1515 920 1519
rect 935 1515 939 1519
rect 910 1397 914 1401
rect 892 1144 896 1148
rect 911 1144 915 1148
rect 838 1069 842 1073
rect 831 1059 835 1063
rect 138 1041 142 1045
rect 207 1041 211 1045
rect 234 1029 238 1033
rect 830 1029 834 1033
rect 140 1010 144 1014
rect 817 999 821 1003
rect -611 967 -607 971
rect 691 968 695 972
rect 926 969 930 973
rect 134 959 138 963
rect 905 959 909 963
rect 921 959 925 963
rect 768 952 773 957
rect 906 952 910 956
rect 925 952 929 956
rect -233 917 -229 921
rect -224 917 -220 921
rect -343 910 -339 914
rect -233 899 -229 903
rect -224 901 -220 905
rect -118 917 -114 921
rect -127 903 -123 907
rect 12 936 16 940
rect 26 936 30 940
rect 145 936 149 940
rect 12 911 16 915
rect 159 936 163 940
rect 817 939 821 943
rect 827 939 831 943
rect 873 932 877 936
rect 270 924 274 928
rect 601 924 605 928
rect 197 917 201 921
rect 26 910 30 914
rect 56 910 60 914
rect 142 910 146 914
rect 169 910 173 914
rect 190 910 194 914
rect 505 910 509 914
rect 135 903 139 907
rect -224 885 -220 889
rect -97 887 -93 891
rect -67 889 -63 893
rect 135 895 139 899
rect -220 858 -216 862
rect 132 887 136 891
rect 12 879 16 883
rect 169 896 173 900
rect 613 909 617 913
rect 622 900 626 904
rect 190 895 194 899
rect 601 886 605 890
rect 817 921 821 925
rect 827 921 831 925
rect 838 923 842 927
rect 873 908 877 912
rect 880 932 884 936
rect 924 932 928 936
rect 917 923 921 927
rect 880 908 884 912
rect 817 901 821 905
rect 827 901 831 905
rect 902 901 906 905
rect 962 1024 966 1028
rect 945 969 949 973
rect 944 960 948 964
rect 943 952 947 956
rect 1640 953 1644 957
rect 952 946 956 950
rect 979 945 983 949
rect 951 939 955 943
rect 1004 938 1008 942
rect 942 932 946 936
rect 978 931 982 935
rect 959 925 963 929
rect 1444 924 1448 928
rect 1383 914 1387 918
rect 989 910 993 914
rect 781 890 785 894
rect 817 887 821 891
rect 146 858 150 862
rect 628 858 632 862
rect 88 853 92 857
rect 88 407 92 411
rect 88 386 92 390
rect 26 289 30 293
rect 860 879 864 883
rect 1472 886 1476 890
rect 994 859 998 863
rect 1476 858 1480 862
rect 937 409 941 413
rect 937 392 941 396
rect 874 289 878 293
rect 842 260 846 264
rect 1680 961 1684 965
rect 1752 960 1756 964
rect 1722 944 1726 948
rect 1752 945 1756 949
rect 1673 935 1677 939
rect 1708 879 1712 883
rect 1722 289 1726 293
rect 1718 268 1722 272
rect 1679 261 1683 265
rect 3 256 7 260
rect 88 256 92 260
rect 937 257 941 261
rect 1792 260 1796 264
rect 1792 244 1796 248
rect 125 181 129 185
rect 89 172 93 176
rect 973 181 977 185
rect 937 172 941 176
<< metal2 >>
rect -761 2620 -751 2623
rect 50 2621 98 2624
rect 896 2620 945 2623
rect 1745 2621 1797 2624
rect -761 1886 -758 2620
rect 101 2528 163 2531
rect -729 2526 -681 2527
rect -742 2524 -681 2526
rect -742 2523 -699 2524
rect -742 1933 -739 2523
rect -731 2513 -701 2517
rect -731 2508 -727 2513
rect -684 2510 -681 2524
rect -693 2507 -681 2510
rect -485 1948 -481 1953
rect -447 1951 -405 1954
rect -485 1944 -455 1948
rect -742 1930 -734 1933
rect -737 1907 -734 1930
rect -697 1911 -678 1914
rect -697 1907 -694 1911
rect -737 1904 -694 1907
rect -681 1907 -678 1911
rect -675 1913 -672 1930
rect -675 1910 -634 1913
rect -681 1904 -647 1907
rect -690 1886 -687 1904
rect -761 1883 -687 1886
rect -650 1854 -647 1904
rect -637 1901 -634 1910
rect -608 1908 -604 1918
rect -577 1908 -574 1919
rect -451 1905 -447 1916
rect -637 1898 -561 1901
rect -624 1858 -571 1862
rect -650 1851 -571 1854
rect -564 1848 -561 1898
rect -408 1873 -405 1951
rect -3 1948 1 1953
rect 35 1951 46 1954
rect -3 1944 27 1948
rect -362 1880 -358 1921
rect -331 1866 -328 1894
rect -36 1873 -33 1884
rect -319 1870 -33 1873
rect 43 1874 46 1951
rect 101 1933 104 2528
rect 117 2513 147 2517
rect 117 2508 121 2513
rect 160 2510 163 2528
rect 155 2507 163 2510
rect 933 2418 937 2515
rect 965 2513 995 2517
rect 965 2508 969 2513
rect 1029 2510 1032 2541
rect 1003 2507 1032 2510
rect 1794 2398 1797 2621
rect 1782 2395 1797 2398
rect 363 1948 367 1953
rect 401 1951 444 1954
rect 363 1944 393 1948
rect 89 1930 105 1933
rect 89 1887 92 1930
rect 117 1896 121 1919
rect 151 1918 157 1921
rect 117 1892 143 1896
rect 89 1884 124 1887
rect 121 1881 124 1884
rect 139 1881 143 1892
rect 154 1881 157 1918
rect 172 1881 175 1930
rect 214 1881 218 1913
rect 240 1897 244 1916
rect 269 1898 272 1919
rect 397 1883 401 1916
rect 441 1887 444 1951
rect 845 1948 849 1953
rect 883 1951 892 1954
rect 889 1948 892 1951
rect 845 1944 875 1948
rect 889 1909 892 1943
rect 933 1927 937 2388
rect 1211 1948 1215 1953
rect 1249 1951 1261 1954
rect 1211 1944 1241 1948
rect 999 1918 1017 1921
rect 895 1914 929 1917
rect 895 1909 898 1914
rect 926 1909 929 1914
rect 945 1911 1037 1914
rect 945 1909 948 1911
rect 889 1906 898 1909
rect 926 1906 948 1909
rect 1034 1909 1037 1911
rect 718 1899 890 1902
rect 502 1887 505 1893
rect 441 1884 505 1887
rect 397 1879 416 1883
rect 517 1874 520 1895
rect 536 1883 539 1893
rect 43 1871 520 1874
rect -331 1863 80 1866
rect 111 1864 128 1868
rect -639 1845 -628 1848
rect -564 1845 67 1848
rect -642 971 -638 1840
rect -631 1684 -628 1845
rect -620 1834 -616 1837
rect -619 1825 -616 1834
rect -619 1822 -590 1825
rect -593 1790 -590 1822
rect 77 1776 80 1863
rect 155 1861 159 1863
rect 111 1858 159 1861
rect 107 1845 125 1848
rect 109 1835 150 1838
rect 109 1826 163 1830
rect 84 1742 88 1782
rect 78 1738 88 1742
rect -633 1680 -628 1684
rect -633 977 -630 1680
rect 138 1410 144 1413
rect 151 1392 154 1817
rect 143 1389 154 1392
rect 76 1301 126 1304
rect 76 1294 80 1301
rect 112 1290 124 1294
rect 83 1260 87 1286
rect 78 1256 87 1260
rect 136 1122 140 1383
rect 143 1305 146 1389
rect 159 1294 163 1826
rect 172 1817 175 1864
rect 718 1840 721 1899
rect 911 1896 915 1905
rect 731 1892 915 1896
rect 731 1850 735 1892
rect 931 1871 932 1875
rect 919 1856 922 1863
rect 928 1864 932 1871
rect 965 1864 969 1904
rect 928 1860 969 1864
rect 1034 1906 1050 1909
rect 1018 1856 1021 1904
rect 843 1852 912 1855
rect 919 1853 1021 1856
rect 731 1849 831 1850
rect 731 1847 888 1849
rect 731 1846 884 1847
rect 909 1847 912 1852
rect 909 1844 1021 1847
rect 1028 1841 1031 1904
rect 1047 1889 1050 1906
rect 1088 1897 1092 1917
rect 1119 1897 1122 1919
rect 1249 1907 1253 1918
rect 1151 1901 1244 1904
rect 1151 1890 1155 1901
rect 1089 1889 1155 1890
rect 1047 1886 1155 1889
rect 1241 1895 1244 1901
rect 1258 1902 1261 1951
rect 1693 1948 1697 1953
rect 1731 1951 1740 1954
rect 1693 1944 1723 1948
rect 1334 1895 1338 1896
rect 1241 1892 1338 1895
rect 1221 1889 1225 1892
rect 1365 1889 1368 1893
rect 1221 1885 1368 1889
rect 1737 1866 1740 1951
rect 1782 1910 1785 2395
rect 1537 1863 1740 1866
rect 1763 1907 1785 1910
rect 1237 1857 1505 1860
rect 1226 1851 1500 1854
rect 718 1837 891 1840
rect 905 1838 1031 1841
rect 905 1831 908 1838
rect 1258 1835 1263 1838
rect 147 1290 163 1294
rect 166 1814 175 1817
rect 863 1828 908 1831
rect 921 1832 1263 1835
rect 1537 1834 1541 1863
rect 166 1188 169 1814
rect 826 1799 830 1826
rect 839 1777 843 1822
rect 236 1773 246 1777
rect 835 1773 843 1777
rect 236 1747 240 1773
rect 832 1743 851 1746
rect 243 1686 246 1740
rect 198 1683 246 1686
rect 198 1627 201 1683
rect 680 1670 683 1684
rect 213 1667 683 1670
rect 693 1664 696 1694
rect 769 1687 772 1693
rect 724 1684 772 1687
rect 863 1667 866 1828
rect 921 1823 925 1832
rect 1388 1831 1541 1834
rect 1560 1855 1690 1859
rect 1712 1856 1751 1859
rect 1388 1829 1391 1831
rect 869 1819 925 1823
rect 929 1826 1391 1829
rect 869 1673 873 1819
rect 929 1816 932 1826
rect 877 1813 932 1816
rect 877 1679 881 1813
rect 888 1796 938 1800
rect 1527 1796 1536 1800
rect 1532 1770 1536 1796
rect 895 1766 937 1769
rect 1560 1766 1564 1855
rect 1570 1849 1683 1852
rect 1526 1756 1529 1762
rect 1570 1756 1573 1849
rect 1639 1820 1642 1840
rect 884 1752 943 1755
rect 1526 1753 1573 1756
rect 884 1688 887 1752
rect 877 1676 894 1679
rect 869 1670 886 1673
rect 863 1664 880 1667
rect 693 1661 849 1664
rect 208 1654 211 1658
rect 798 1654 807 1658
rect 803 1628 807 1654
rect 198 1624 211 1627
rect 846 1625 849 1661
rect 270 1545 273 1574
rect 187 1542 273 1545
rect 347 1545 350 1574
rect 797 1569 800 1620
rect 797 1566 846 1569
rect 347 1542 867 1545
rect 187 1442 190 1542
rect 236 1535 246 1539
rect 236 1509 240 1535
rect 243 1454 246 1501
rect 197 1451 246 1454
rect 187 1439 217 1442
rect 682 1426 685 1446
rect 172 1423 685 1426
rect 694 1427 697 1456
rect 769 1449 772 1455
rect 721 1446 772 1449
rect 694 1424 831 1427
rect 172 1336 175 1423
rect 798 1416 807 1420
rect 803 1390 807 1416
rect 797 1353 800 1382
rect 828 1360 831 1424
rect 828 1357 857 1360
rect 797 1350 854 1353
rect 172 1333 193 1336
rect 190 1323 193 1333
rect 271 1331 274 1336
rect 255 1328 274 1331
rect 346 1316 349 1336
rect 178 1313 349 1316
rect 236 1297 245 1301
rect 835 1297 841 1301
rect 180 1280 189 1283
rect 236 1271 240 1297
rect 851 1270 854 1350
rect 832 1267 854 1270
rect 243 1223 246 1263
rect 864 1243 867 1542
rect 823 1240 867 1243
rect 194 1220 246 1223
rect 673 1188 676 1208
rect 166 1185 676 1188
rect 693 1190 696 1217
rect 770 1211 773 1217
rect 705 1208 773 1211
rect 877 1190 880 1664
rect 883 1637 886 1670
rect 890 1431 894 1676
rect 907 1673 936 1677
rect 934 1646 937 1647
rect 926 1643 937 1646
rect 926 1636 929 1643
rect 905 1633 929 1636
rect 964 1550 974 1554
rect 963 1524 967 1550
rect 905 1515 916 1519
rect 920 1515 935 1519
rect 972 1504 975 1516
rect 903 1501 975 1504
rect 890 1427 915 1431
rect 693 1187 880 1190
rect 796 1178 805 1182
rect 147 1164 172 1167
rect 147 1133 158 1137
rect 118 1118 140 1122
rect -539 1052 -476 1055
rect -539 977 -536 1052
rect -479 1048 -476 1052
rect -486 1014 -482 1040
rect -486 1010 -476 1014
rect -633 974 -536 977
rect 118 976 122 1118
rect 169 1110 172 1164
rect 177 1143 180 1178
rect 801 1152 805 1178
rect 177 1140 212 1143
rect 149 1107 172 1110
rect 129 1070 139 1073
rect 129 1041 138 1044
rect 129 1010 140 1014
rect -86 971 122 976
rect -642 967 -611 971
rect -86 962 -82 971
rect -233 958 -82 962
rect 12 959 134 962
rect -233 921 -230 958
rect 12 940 15 959
rect 149 954 153 1107
rect 176 1102 180 1133
rect 209 1122 212 1140
rect 209 1119 218 1122
rect 795 1104 798 1144
rect 157 1098 180 1102
rect 157 961 161 1098
rect 268 1091 271 1099
rect 268 1088 326 1091
rect 345 1070 348 1103
rect 795 1101 855 1104
rect 818 1088 841 1091
rect 358 1076 361 1088
rect 811 1076 814 1088
rect 358 1073 814 1076
rect 818 1070 821 1088
rect 345 1067 821 1070
rect 838 1073 841 1088
rect 845 1063 849 1094
rect 234 1059 244 1063
rect 835 1059 849 1063
rect 211 1041 213 1045
rect 210 1018 213 1041
rect 234 1033 238 1059
rect 852 1032 855 1101
rect 834 1029 855 1032
rect 241 1018 244 1029
rect 210 1015 244 1018
rect 858 1003 861 1174
rect 892 1148 896 1401
rect 900 1141 903 1420
rect 915 1144 947 1148
rect 900 1138 930 1141
rect 927 1038 930 1138
rect 821 1000 861 1003
rect 915 1035 930 1038
rect 691 972 694 979
rect 157 957 194 961
rect 149 951 172 954
rect 149 936 159 939
rect -92 929 146 933
rect -220 917 -118 921
rect -92 914 -88 929
rect -313 912 -88 914
rect -310 910 -88 912
rect -84 920 113 923
rect -84 906 -81 920
rect -123 903 -81 906
rect -233 855 -230 899
rect -224 889 -220 901
rect 12 883 15 911
rect 26 885 29 910
rect 56 888 60 910
rect 110 884 113 920
rect 142 914 146 929
rect 169 914 172 951
rect 190 914 194 957
rect 768 957 771 979
rect 874 959 905 962
rect 793 948 842 952
rect 206 944 796 948
rect 206 920 210 944
rect 535 931 714 935
rect 201 917 210 920
rect 270 907 274 924
rect 535 913 539 931
rect 139 903 274 907
rect 139 896 169 899
rect 190 891 194 895
rect 136 887 194 891
rect 601 890 605 924
rect 711 914 714 931
rect 817 925 821 939
rect 827 925 830 939
rect 838 927 842 948
rect 874 936 877 959
rect 880 952 906 956
rect 880 936 884 952
rect 915 942 918 1035
rect 943 1031 947 1144
rect 962 1068 972 1072
rect 943 1028 956 1031
rect 930 969 945 972
rect 925 960 944 963
rect 929 952 943 956
rect 952 950 956 1028
rect 962 1028 966 1068
rect 915 939 951 942
rect 928 932 942 936
rect 852 925 911 929
rect 852 920 855 925
rect 842 918 855 920
rect 751 917 855 918
rect 858 917 903 921
rect 751 914 846 917
rect 617 909 695 912
rect 711 910 754 914
rect 858 913 861 917
rect 850 911 861 913
rect 900 913 903 917
rect 907 920 911 925
rect 921 924 959 928
rect 969 928 972 1037
rect 1680 965 1683 1849
rect 1686 972 1690 1855
rect 1705 1850 1751 1853
rect 1763 1843 1766 1907
rect 1719 1840 1766 1843
rect 1686 968 1756 972
rect 1752 964 1756 968
rect 1644 953 1789 957
rect 983 945 1633 949
rect 1008 939 1602 942
rect 982 931 1476 935
rect 969 924 1011 928
rect 907 916 993 920
rect 989 914 993 916
rect 1008 917 1011 924
rect 1008 914 1356 917
rect 762 910 861 911
rect 613 908 695 909
rect 691 904 695 908
rect 762 908 853 910
rect 762 904 765 908
rect 691 901 765 904
rect 622 891 625 900
rect 616 887 625 891
rect 817 891 820 901
rect 827 896 830 901
rect 827 893 839 896
rect 836 891 839 893
rect 836 888 863 891
rect 110 881 136 884
rect -216 858 -186 862
rect -233 852 -224 855
rect -190 853 -186 858
rect 88 411 92 853
rect 133 855 136 881
rect 150 858 180 861
rect 133 852 142 855
rect 176 853 179 858
rect 616 855 619 887
rect 860 883 863 888
rect 874 885 877 908
rect 900 910 964 913
rect 1353 911 1356 914
rect 880 895 884 908
rect 906 901 955 905
rect 880 891 908 895
rect 904 888 908 891
rect 632 858 662 862
rect 616 852 624 855
rect 658 853 662 858
rect 951 784 955 901
rect 961 856 964 910
rect 998 859 1027 862
rect 1006 858 1027 859
rect 961 853 993 856
rect 1024 853 1027 858
rect 1444 855 1447 924
rect 1472 890 1476 931
rect 1598 887 1602 939
rect 1629 888 1633 945
rect 1677 935 1711 938
rect 1708 883 1711 935
rect 1722 885 1725 944
rect 1752 888 1756 945
rect 1480 858 1510 862
rect 1444 852 1475 855
rect 1506 853 1510 858
rect 938 780 955 784
rect 938 413 942 780
rect 941 409 942 413
rect 3 297 23 300
rect 3 260 6 297
rect 56 293 60 299
rect 30 289 60 293
rect 88 260 92 386
rect 842 296 871 299
rect 842 264 846 296
rect 904 293 908 299
rect 878 289 908 293
rect 937 261 941 392
rect 1679 296 1719 299
rect 1679 265 1682 296
rect 1752 293 1756 298
rect 1726 289 1756 293
rect 1785 272 1789 953
rect 1722 268 1789 272
rect 1792 248 1795 260
rect 79 186 128 189
rect 927 186 976 189
rect 125 185 128 186
rect 973 185 976 186
rect 89 155 93 172
rect 937 155 941 172
<< m1p >>
rect 910 1397 914 1401
use top_bott_tree  top_bott_tree_1
timestamp 1383892968
transform -1 0 1016 0 -1 2799
box -775 129 1777 907
use new_tree  new_tree_0
timestamp 1383892968
transform 0 1 -516 -1 0 1828
box -8 -123 848 655
use lut  lut_6
timestamp 1383712281
transform 1 0 242 0 1 1693
box -34 0 593 108
use lut  lut_5
timestamp 1383712281
transform -1 0 801 0 1 1574
box -34 0 593 108
use lut  lut_4
timestamp 1383712281
transform 1 0 242 0 1 1455
box -34 0 593 108
use lut  lut_3
timestamp 1383712281
transform -1 0 801 0 1 1336
box -34 0 593 108
use lut  lut_2
timestamp 1383712281
transform 1 0 242 0 1 1217
box -34 0 593 108
use lut  lut_1
timestamp 1383712281
transform -1 0 799 0 1 1098
box -34 0 593 108
use lut  lut_0
timestamp 1383712281
transform 1 0 240 0 1 979
box -34 0 593 108
use new_tree  new_tree_1
timestamp 1383892968
transform 0 -1 1566 1 0 982
box -8 -123 848 655
use mux  mux_0
timestamp 1382957000
transform 1 0 -772 0 1 897
box -2 0 71 108
use mux  mux_1
timestamp 1382957000
transform 1 0 -712 0 1 897
box -2 0 71 108
use top_bott_tree  top_bott_tree_0
timestamp 1383892968
transform 1 0 9 0 1 7
box -775 129 1777 907
<< end >>
