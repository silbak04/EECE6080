magic
tech scmos
timestamp 1383633248
<< error_s >>
rect -524 586 -521 590
<< metal1 >>
rect -755 1020 -739 1023
rect 74 615 87 616
rect 74 613 90 615
rect 97 614 99 615
rect -761 587 -525 590
rect -761 552 -525 555
rect 67 507 70 575
rect 74 532 77 613
rect 87 609 90 613
rect 98 612 99 614
rect 98 603 108 606
rect 94 593 97 595
rect 87 569 90 590
rect 94 569 97 572
rect 87 531 90 550
rect 94 532 97 550
rect 87 520 90 528
rect 87 516 88 520
rect 87 507 90 516
rect 67 504 87 507
rect -755 499 -701 502
rect -97 499 -80 502
rect -755 490 -701 493
rect -747 -33 -737 -30
rect -738 -34 -737 -33
rect -747 -123 -738 -120
rect -816 -133 -807 -130
rect -816 -188 -807 -185
rect -816 -196 -807 -193
rect -816 -204 -807 -201
<< m2contact >>
rect -759 1019 -755 1023
rect -739 1019 -735 1023
rect -765 587 -761 591
rect -525 586 -521 590
rect 67 575 71 579
rect -765 552 -761 556
rect 128 611 132 615
rect 74 528 78 532
rect -759 499 -755 503
rect -701 499 -697 503
rect -101 498 -97 502
rect -80 498 -76 502
rect -759 490 -755 494
rect -701 490 -697 494
rect -751 -34 -747 -30
rect -722 -44 -718 -40
rect -751 -123 -747 -119
rect -630 -120 -626 -116
rect -820 -134 -816 -130
rect -807 -134 -803 -130
rect -720 -134 -716 -130
rect -696 -134 -692 -130
rect -688 -134 -684 -130
rect -680 -134 -676 -130
rect -672 -134 -668 -130
rect -648 -134 -644 -130
rect -820 -189 -816 -185
rect -807 -189 -803 -185
rect -820 -197 -816 -193
rect -807 -197 -803 -193
rect -820 -205 -816 -201
rect -807 -205 -803 -201
<< metal2 >>
rect -819 1287 79 1290
rect -819 -130 -816 1287
rect -813 1263 87 1266
rect -813 -208 -810 1263
rect -807 1122 -641 1125
rect -807 83 -804 1122
rect -801 1112 -640 1115
rect -801 117 -798 1112
rect -795 1071 -711 1074
rect -795 195 -792 1071
rect -789 1065 -712 1068
rect -789 230 -786 1065
rect -783 1059 -712 1062
rect -783 264 -780 1059
rect -777 1053 -704 1056
rect -777 270 -774 1053
rect -771 1047 -711 1050
rect -771 555 -768 1047
rect -765 1041 -710 1044
rect -765 591 -762 1041
rect -752 1032 -711 1035
rect -771 552 -765 555
rect -758 503 -755 1019
rect -758 276 -755 490
rect -752 285 -749 1032
rect -746 1026 -712 1029
rect -746 291 -743 1026
rect -735 1020 -696 1023
rect -740 985 -708 988
rect -740 297 -737 985
rect -734 951 -708 954
rect -734 303 -731 951
rect -728 872 -708 875
rect -728 309 -725 872
rect -722 838 -709 841
rect -722 315 -719 838
rect -716 760 -708 763
rect -716 357 -713 760
rect -709 388 -706 725
rect 46 609 63 612
rect 51 587 57 590
rect 54 559 57 587
rect 60 569 63 609
rect 129 579 132 611
rect 71 576 132 579
rect 60 566 1761 569
rect 54 556 1761 559
rect 48 550 51 556
rect 48 547 1761 550
rect -697 499 -101 502
rect -91 493 -87 506
rect -15 502 -11 506
rect -76 499 -11 502
rect -697 490 -87 493
rect -709 385 -639 388
rect -716 354 -642 357
rect -722 312 -711 315
rect -728 306 -712 309
rect -734 300 -710 303
rect -740 294 -712 297
rect -746 288 -709 291
rect -752 282 -711 285
rect -758 273 -712 276
rect -777 267 -708 270
rect -783 261 -690 264
rect -789 227 -708 230
rect -795 192 -709 195
rect -801 114 -703 117
rect -807 80 -709 83
rect -722 0 -708 4
rect -751 -119 -748 -34
rect -722 -40 -719 0
rect -709 -77 -706 -34
rect -709 -80 -627 -77
rect -630 -116 -627 -80
rect -803 -133 -720 -130
rect -696 -186 -693 -134
rect -803 -189 -693 -186
rect -684 -194 -680 -130
rect -803 -197 -680 -194
rect -672 -202 -669 -134
rect -803 -205 -669 -202
rect -648 -208 -645 -134
rect -813 -211 -645 -208
use lut  lut_1
timestamp 1383530834
transform 1 0 -600 0 1 1408
box 0 0 593 108
use shift_slice  shift_slice_0
timestamp 1383130333
transform 1 0 953 0 1 1421
box 0 0 112 108
use lut_p_tree  lut_p_tree_1
timestamp 1383633248
transform 1 0 -630 0 1 576
box -82 -10 2429 733
use lut  lut_0
timestamp 1383530834
transform 1 0 -542 0 1 506
box 0 0 593 108
use BUFX4  BUFX4_0
timestamp 1053722803
transform 1 0 -740 0 1 -77
box -9 -3 37 105
use mux  mux_0
timestamp 1382957000
transform -1 0 -679 0 -1 -84
box -2 0 71 108
use mux  mux_1
timestamp 1382957000
transform 1 0 -685 0 -1 -84
box -2 0 71 108
use lut_p_tree  lut_p_tree_0
timestamp 1383633248
transform 1 0 -630 0 1 -183
box -82 -10 2429 733
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 -368 0 1 -486
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_0
timestamp 1383129201
transform 1 0 -76 0 1 -483
box -8 -3 104 105
<< end >>
