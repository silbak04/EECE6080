magic
tech scmos
timestamp 1384231894
<< error_s >>
rect 3 8 4 10
<< metal1 >>
rect 2 100 6 106
rect 7 45 21 48
rect 102 46 105 50
rect 8 36 14 39
rect 103 0 109 6
use DFFPOSX1  DFFPOSX1_0
timestamp 1384231894
transform 1 0 8 0 1 3
box -8 -5 104 105
<< labels >>
rlabel metal1 3 103 3 103 6 VDD
rlabel metal1 8 46 8 46 6 P_IN
rlabel metal1 9 37 9 37 6 PCLKI
rlabel metal1 104 48 104 48 6 P_OUT
rlabel metal1 104 3 104 3 6 GND
<< end >>
