magic
tech scmos
timestamp 1383648289
<< error_s >>
rect -524 586 -521 590
<< metal1 >>
rect -840 1316 1820 1325
rect -840 1309 -832 1316
rect -840 1306 83 1309
rect -840 1303 86 1306
rect -840 1196 -832 1303
rect 1812 1196 1820 1312
rect -840 1190 -642 1196
rect 1744 1190 1820 1196
rect -840 911 -832 1190
rect -822 1090 -642 1096
rect 1744 1090 1803 1096
rect 1812 1083 1820 1190
rect 1744 1077 1820 1083
rect -119 1032 -90 1038
rect -755 1020 -739 1023
rect -822 1005 -711 1011
rect -119 1005 -113 1032
rect 1744 977 1803 983
rect 1812 970 1820 1077
rect 1744 964 1820 970
rect -840 905 -706 911
rect -840 798 -832 905
rect -822 892 -711 898
rect 1744 864 1803 870
rect -840 792 -706 798
rect -840 685 -832 792
rect -822 779 -711 785
rect 1642 779 1803 785
rect 1812 685 1820 964
rect -840 679 -706 685
rect 1642 679 1820 685
rect -840 512 -832 679
rect 917 666 1803 672
rect 74 615 87 616
rect 74 613 90 615
rect 97 614 99 615
rect -822 606 -541 612
rect -761 587 -525 590
rect -761 552 -525 555
rect -840 506 -536 512
rect 67 507 70 575
rect 74 532 77 613
rect 87 609 90 613
rect 98 612 99 614
rect 98 603 108 606
rect 94 593 97 595
rect 87 569 90 590
rect 1812 572 1820 679
rect 94 569 97 572
rect 917 566 1820 572
rect 1812 550 1820 566
rect 87 531 90 550
rect 94 532 97 550
rect 918 544 1820 550
rect 87 520 90 528
rect 87 516 88 520
rect 87 507 90 516
rect -840 152 -832 506
rect 67 504 87 507
rect -755 499 -701 502
rect -97 499 -80 502
rect -755 490 -701 493
rect 918 444 1803 450
rect 1812 437 1820 544
rect 1744 431 1820 437
rect 1744 331 1803 337
rect 1812 324 1820 431
rect 1744 318 1820 324
rect -125 273 -90 279
rect -125 252 -119 273
rect -823 246 -711 252
rect 1744 218 1803 224
rect 1812 211 1820 318
rect 1744 205 1820 211
rect -840 146 -706 152
rect -840 39 -832 146
rect -823 133 -711 139
rect 1744 105 1803 111
rect -840 33 -706 39
rect -840 -74 -832 33
rect -823 20 -742 26
rect 1642 20 1803 26
rect -747 -33 -737 -30
rect -738 -34 -737 -33
rect 1812 -74 1820 205
rect -840 -80 -740 -74
rect 1642 -80 1820 -74
rect -840 -84 -832 -80
rect -840 -90 -741 -84
rect -840 -216 -832 -90
rect 917 -93 1803 -87
rect -747 -123 -738 -120
rect -816 -133 -807 -130
rect -823 -179 -756 -173
rect -763 -184 -756 -179
rect -816 -188 -807 -185
rect -763 -190 -740 -184
rect 1812 -187 1820 -80
rect 917 -193 1820 -187
rect -816 -196 -807 -193
rect -816 -204 -807 -201
rect 1812 -216 1820 -193
rect -840 -224 1820 -216
<< m2contact >>
rect -850 1090 -843 1096
rect -849 1005 -843 1011
rect -829 1090 -822 1096
rect 1803 1090 1809 1096
rect 1823 1090 1829 1096
rect -759 1019 -755 1023
rect -739 1019 -735 1023
rect -828 1005 -822 1011
rect 1803 977 1809 983
rect 1823 977 1829 983
rect -849 892 -843 898
rect -828 892 -822 898
rect 1803 864 1809 870
rect -849 779 -843 785
rect -828 779 -822 785
rect 1803 779 1809 785
rect 1823 864 1829 870
rect 1823 779 1829 785
rect -850 606 -844 612
rect 1803 666 1809 672
rect -828 606 -822 612
rect -765 587 -761 591
rect -525 586 -521 590
rect 67 575 71 579
rect -765 552 -761 556
rect 128 611 132 615
rect 1823 666 1829 672
rect 74 528 78 532
rect -849 246 -843 252
rect -759 499 -755 503
rect -701 499 -697 503
rect -101 498 -97 502
rect -80 498 -76 502
rect -759 490 -755 494
rect -701 490 -697 494
rect 1803 444 1809 450
rect 1823 444 1829 450
rect 1803 331 1809 337
rect 1823 331 1829 337
rect -829 246 -823 252
rect 1803 218 1809 224
rect 1823 218 1829 224
rect -849 133 -843 139
rect -829 133 -823 139
rect 1803 105 1809 111
rect -849 20 -843 26
rect -829 20 -823 26
rect 1803 20 1809 26
rect -751 -34 -747 -30
rect -722 -44 -718 -40
rect 1823 105 1829 111
rect 1823 20 1829 26
rect -849 -179 -843 -173
rect 1803 -93 1809 -87
rect -751 -123 -747 -119
rect -630 -120 -626 -116
rect -820 -134 -816 -130
rect -807 -134 -803 -130
rect -720 -134 -716 -130
rect -696 -134 -692 -130
rect -688 -134 -684 -130
rect -680 -134 -676 -130
rect -672 -134 -668 -130
rect -648 -134 -644 -130
rect -829 -179 -823 -173
rect -820 -189 -816 -185
rect -807 -189 -803 -185
rect 1823 -93 1829 -87
rect -820 -197 -816 -193
rect -807 -197 -803 -193
rect -820 -205 -816 -201
rect -807 -205 -803 -201
<< metal2 >>
rect -819 1287 79 1290
rect -843 1090 -829 1096
rect -843 1005 -828 1011
rect -843 892 -828 898
rect -843 779 -828 785
rect -844 606 -828 612
rect -843 246 -829 252
rect -843 133 -829 139
rect -843 20 -829 26
rect -819 -130 -816 1287
rect -813 1263 87 1266
rect -843 -179 -829 -173
rect -813 -208 -810 1263
rect -807 1122 -641 1125
rect -807 83 -804 1122
rect -801 1112 -640 1115
rect -801 117 -798 1112
rect 1809 1090 1823 1096
rect -795 1071 -711 1074
rect -795 195 -792 1071
rect -789 1065 -712 1068
rect -789 230 -786 1065
rect -783 1059 -712 1062
rect -783 264 -780 1059
rect -777 1053 -704 1056
rect -777 270 -774 1053
rect -771 1047 -711 1050
rect -771 555 -768 1047
rect -765 1041 -710 1044
rect -765 591 -762 1041
rect -752 1032 -711 1035
rect -771 552 -765 555
rect -758 503 -755 1019
rect -758 276 -755 490
rect -752 285 -749 1032
rect -746 1026 -712 1029
rect -746 291 -743 1026
rect -735 1020 -696 1023
rect -740 985 -708 988
rect -740 297 -737 985
rect 1809 977 1823 983
rect -734 951 -708 954
rect -734 303 -731 951
rect -728 872 -708 875
rect -728 309 -725 872
rect 1809 864 1823 870
rect -722 838 -709 841
rect -722 315 -719 838
rect 1809 779 1823 785
rect -716 760 -708 763
rect -716 357 -713 760
rect -709 388 -706 725
rect 1809 666 1823 672
rect 46 609 63 612
rect 51 587 57 590
rect 54 559 57 587
rect 60 569 63 609
rect 129 579 132 611
rect 71 576 132 579
rect 60 566 1812 569
rect 54 556 1812 559
rect 48 550 51 556
rect 48 547 1812 550
rect -697 499 -101 502
rect -91 493 -87 506
rect -15 502 -11 506
rect -76 499 -11 502
rect -697 490 -87 493
rect 1809 444 1823 450
rect -709 385 -639 388
rect -716 354 -642 357
rect 1809 331 1823 337
rect -722 312 -711 315
rect -728 306 -712 309
rect -734 300 -710 303
rect -740 294 -712 297
rect -746 288 -709 291
rect -752 282 -711 285
rect -758 273 -712 276
rect -777 267 -708 270
rect -783 261 -690 264
rect -789 227 -708 230
rect 1809 218 1823 224
rect -795 192 -709 195
rect -801 114 -703 117
rect 1809 105 1823 111
rect -807 80 -709 83
rect 1809 20 1823 26
rect -722 0 -708 4
rect -751 -119 -748 -34
rect -722 -40 -719 0
rect -709 -77 -706 -34
rect -709 -80 -627 -77
rect -630 -116 -627 -80
rect 1809 -93 1823 -87
rect -803 -133 -720 -130
rect -696 -186 -693 -134
rect -803 -189 -693 -186
rect -684 -194 -680 -130
rect -803 -197 -680 -194
rect -672 -202 -669 -134
rect -803 -205 -669 -202
rect -648 -208 -645 -134
rect -813 -211 -645 -208
use lut_p_tree  lut_p_tree_1
timestamp 1383647959
transform 1 0 -630 0 1 576
box -82 -10 2429 733
use lut  lut_0
timestamp 1383530834
transform 1 0 -542 0 1 506
box 0 0 593 108
use BUFX4  BUFX4_0
timestamp 1053722803
transform 1 0 -740 0 1 -77
box -9 -3 37 105
use mux  mux_0
timestamp 1382957000
transform -1 0 -679 0 -1 -84
box -2 0 71 108
use mux  mux_1
timestamp 1382957000
transform 1 0 -685 0 -1 -84
box -2 0 71 108
use lut_p_tree  lut_p_tree_0
timestamp 1383647959
transform 1 0 -630 0 1 -183
box -82 -10 2429 733
<< end >>
