magic
tech scmos
timestamp 1384225954
<< metal2 >>
rect 1023 4743 1277 4997
rect 1323 4743 1577 4997
rect 1623 4743 1877 4997
rect 1923 4743 2177 4997
rect 2223 4743 2477 4997
rect 2523 4743 2777 4997
rect 2823 4743 3077 4997
rect 3123 4743 3377 4997
rect 3423 4743 3677 4997
rect 3723 4743 3977 4997
rect 3 3123 257 3377
rect 4743 3123 4997 3377
rect 3 2823 257 3077
rect 4743 2823 4997 3077
rect 3 2523 257 2777
rect 4743 2523 4997 2777
rect 3 2223 257 2477
rect 4743 2223 4997 2477
rect 3 1923 257 2177
rect 4743 1923 4997 2177
rect 3 1623 257 1877
rect 4743 1623 4997 1877
rect 1023 3 1277 257
rect 1323 3 1577 257
rect 1623 3 1877 257
rect 1923 3 2177 257
rect 2223 3 2477 257
rect 2523 3 2777 257
rect 2823 3 3077 257
rect 3123 3 3377 257
rect 3423 3 3677 257
use top  top_0
timestamp 1384219646
transform 1 0 3182 0 1 2064
box -3182 -2064 1818 2936
<< labels >>
rlabel metal2 3 3123 257 3377 0 LO_4
rlabel metal2 3 2823 257 3077 0 PCLKI
rlabel metal2 3 2523 257 2777 0 LCLKI
rlabel metal2 3 2223 257 2477 0 P_IN
rlabel metal2 3 1923 257 2177 0 L_IN
rlabel metal2 3 1623 257 1877 0 TMEI
rlabel metal2 1023 3 1277 257 0 TII
rlabel metal2 1323 3 1577 257 0 TIO
rlabel metal2 1623 3 1877 257 0 TFDI
rlabel metal2 2223 3 2477 257 0 TPCO
rlabel metal2 2823 3 3077 257 0 TFQO
rlabel metal2 3123 3 3377 257 0 PO_1
rlabel metal2 3423 3 3677 257 0 LO_1
rlabel metal2 4743 1623 4997 1877 0 TEMO
rlabel metal2 4743 1923 4997 2177 0 L_OUT
rlabel metal2 4743 2223 4997 2477 0 P_OUT
rlabel metal2 4743 2523 4997 2777 0 LCLKO
rlabel metal2 4743 2823 4997 3077 0 PCLKO
rlabel metal2 4743 3123 4997 3377 0 F
rlabel metal2 3723 4743 3977 4997 0 TSPO
rlabel metal2 3423 4743 3677 4997 0 TSPI
rlabel metal2 3123 4743 3377 4997 0 TSF
rlabel metal2 2823 4743 3077 4997 0 TSLO
rlabel metal2 2523 4743 2777 4997 0 TSB
rlabel metal2 2223 4743 2477 4997 0 VDD
rlabel metal2 1923 4743 2177 4997 0 TSA
rlabel metal2 1623 4743 1877 4997 0 TSLI
rlabel metal2 1323 4743 1577 4997 0 TSCO
rlabel metal2 1023 4743 1277 4997 0 TSCI
rlabel metal2 1923 3 2177 257 0 TFCI
rlabel metal2 2523 3 2777 257 0 GND
<< end >>
