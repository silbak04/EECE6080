magic
tech scmos
timestamp 1383723055
<< error_s >>
rect 1354 2104 1357 2108
use shift_slice  shift_slice_0
timestamp 1383130333
transform -1 0 1330 0 -1 2307
box 0 0 112 108
use box  box_0
timestamp 1383723055
transform 1 0 1992 0 1 1102
box -770 136 1791 2670
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1072203966
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< end >>
