magic
tech scmos
timestamp 1384231894
<< polysilicon >>
rect 0 0 150 2900
<< end >>
