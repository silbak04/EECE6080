magic
tech scmos
timestamp 1382955972
<< nwell >>
rect 317 427 351 484
rect 420 427 478 484
rect 431 423 458 427
rect 429 294 464 351
rect 416 175 474 232
rect 427 171 454 175
<< ntransistor >>
rect 333 385 335 395
rect 432 389 434 399
rect 440 389 442 409
rect 445 389 447 409
rect 453 389 455 409
rect 458 389 460 409
rect 445 252 447 262
rect 428 137 430 147
rect 436 137 438 157
rect 441 137 443 157
rect 449 137 451 157
rect 454 137 456 157
<< ptransistor >>
rect 333 453 335 473
rect 432 449 434 469
rect 440 429 442 469
rect 445 429 447 469
rect 453 433 455 473
rect 458 433 460 473
rect 445 320 447 340
rect 428 197 430 217
rect 436 177 438 217
rect 441 177 443 217
rect 449 181 451 221
rect 454 181 456 221
<< ndiffusion >>
rect 437 407 440 409
rect 328 394 333 395
rect 332 385 333 394
rect 335 394 340 395
rect 335 385 336 394
rect 431 389 432 399
rect 434 389 435 399
rect 439 389 440 407
rect 442 389 445 409
rect 447 407 453 409
rect 447 389 448 407
rect 452 389 453 407
rect 455 389 458 409
rect 460 389 461 409
rect 440 261 445 262
rect 444 252 445 261
rect 447 261 452 262
rect 447 252 448 261
rect 433 155 436 157
rect 427 137 428 147
rect 430 137 431 147
rect 435 137 436 155
rect 438 137 441 157
rect 443 155 449 157
rect 443 137 444 155
rect 448 137 449 155
rect 451 137 454 157
rect 456 137 457 157
<< pdiffusion >>
rect 328 472 333 473
rect 332 453 333 472
rect 335 472 340 473
rect 335 453 336 472
rect 431 449 432 469
rect 434 449 435 469
rect 439 435 440 469
rect 437 429 440 435
rect 442 429 445 469
rect 447 435 448 469
rect 452 435 453 473
rect 447 433 453 435
rect 455 433 458 473
rect 460 433 461 473
rect 447 429 450 433
rect 440 339 445 340
rect 444 320 445 339
rect 447 339 452 340
rect 447 320 448 339
rect 427 197 428 217
rect 430 197 431 217
rect 435 183 436 217
rect 433 177 436 183
rect 438 177 441 217
rect 443 183 444 217
rect 448 183 449 221
rect 443 181 449 183
rect 451 181 454 221
rect 456 181 457 221
rect 443 177 446 181
<< ndcontact >>
rect 328 385 332 394
rect 336 385 340 394
rect 427 389 431 399
rect 435 389 439 407
rect 448 389 452 407
rect 461 389 465 409
rect 440 252 444 261
rect 448 252 452 261
rect 423 137 427 147
rect 431 137 435 155
rect 444 137 448 155
rect 457 137 461 157
<< pdcontact >>
rect 328 453 332 472
rect 336 453 340 472
rect 427 449 431 469
rect 435 435 439 469
rect 448 435 452 473
rect 461 433 465 473
rect 440 320 444 339
rect 448 320 452 339
rect 423 197 427 217
rect 431 183 435 217
rect 444 183 448 221
rect 457 181 461 221
<< psubstratepcontact >>
rect 324 377 328 381
rect 423 377 427 381
rect 439 377 443 381
rect 455 377 459 381
rect 436 244 440 248
rect 419 125 423 129
rect 435 125 439 129
rect 451 125 455 129
<< nsubstratencontact >>
rect 324 477 328 481
rect 423 477 427 481
rect 439 477 443 481
rect 455 477 459 481
rect 436 344 440 348
rect 419 225 423 229
rect 435 225 439 229
rect 451 225 455 229
<< polysilicon >>
rect 333 473 335 475
rect 432 474 447 476
rect 432 469 434 474
rect 440 469 442 471
rect 445 469 447 474
rect 453 473 455 475
rect 458 473 460 475
rect 333 402 335 453
rect 432 448 434 449
rect 429 446 434 448
rect 429 422 431 446
rect 440 428 442 429
rect 437 426 442 428
rect 445 427 447 429
rect 437 422 439 426
rect 453 419 455 433
rect 458 432 460 433
rect 458 430 461 432
rect 332 398 335 402
rect 429 402 431 418
rect 436 412 438 418
rect 450 417 455 419
rect 445 413 449 415
rect 436 410 442 412
rect 440 409 442 410
rect 445 409 447 413
rect 459 412 461 426
rect 453 409 455 411
rect 458 410 461 412
rect 458 409 460 410
rect 429 400 434 402
rect 432 399 434 400
rect 333 395 335 398
rect 333 383 335 385
rect 432 384 434 389
rect 440 387 442 389
rect 445 387 447 389
rect 453 384 455 389
rect 458 387 460 389
rect 432 382 455 384
rect 445 340 447 342
rect 445 269 447 320
rect 444 265 447 269
rect 445 262 447 265
rect 445 250 447 252
rect 428 222 443 224
rect 428 217 430 222
rect 436 217 438 219
rect 441 217 443 222
rect 449 221 451 223
rect 454 221 456 223
rect 428 196 430 197
rect 425 194 430 196
rect 425 170 427 194
rect 436 176 438 177
rect 433 174 438 176
rect 441 175 443 177
rect 433 170 435 174
rect 449 167 451 181
rect 454 180 456 181
rect 454 178 457 180
rect 425 150 427 166
rect 432 160 434 166
rect 446 165 451 167
rect 441 161 445 163
rect 432 158 438 160
rect 436 157 438 158
rect 441 157 443 161
rect 455 160 457 174
rect 449 157 451 159
rect 454 158 457 160
rect 454 157 456 158
rect 425 148 430 150
rect 428 147 430 148
rect 428 132 430 137
rect 436 135 438 137
rect 441 135 443 137
rect 449 132 451 137
rect 454 135 456 137
rect 428 130 451 132
<< polycontact >>
rect 427 418 431 422
rect 435 418 439 422
rect 328 398 332 402
rect 446 415 450 419
rect 459 426 463 430
rect 440 265 444 269
rect 423 166 427 170
rect 431 166 435 170
rect 442 163 446 167
rect 455 174 459 178
<< metal1 >>
rect 324 481 344 482
rect 328 477 344 481
rect 324 476 344 477
rect 423 481 475 482
rect 427 477 439 481
rect 443 477 455 481
rect 459 477 475 481
rect 423 476 475 477
rect 328 472 332 476
rect 336 472 340 473
rect 435 469 439 476
rect 461 473 465 476
rect 336 420 340 453
rect 427 432 430 449
rect 452 435 456 438
rect 427 430 446 432
rect 328 402 332 406
rect 328 394 332 395
rect 336 394 340 416
rect 427 429 435 430
rect 439 429 446 430
rect 328 382 332 385
rect 324 381 344 382
rect 328 377 344 381
rect 324 376 344 377
rect 203 174 258 178
rect 121 49 125 174
rect 135 166 167 170
rect 254 49 258 174
rect 370 164 374 426
rect 415 422 431 426
rect 377 412 408 416
rect 377 410 381 412
rect 415 371 419 422
rect 435 422 439 426
rect 443 415 446 429
rect 453 416 456 435
rect 463 426 490 430
rect 459 422 463 426
rect 443 413 448 415
rect 427 410 448 413
rect 457 412 463 416
rect 427 399 430 410
rect 453 409 456 412
rect 452 404 456 409
rect 435 382 439 389
rect 461 382 465 389
rect 423 381 475 382
rect 427 377 439 381
rect 443 377 455 381
rect 459 377 475 381
rect 423 376 475 377
rect 415 367 478 371
rect 436 348 456 349
rect 440 344 456 348
rect 436 343 456 344
rect 440 339 444 343
rect 448 339 452 340
rect 448 283 452 320
rect 486 283 490 426
rect 448 279 490 283
rect 440 269 444 273
rect 440 261 444 262
rect 448 261 452 279
rect 440 249 444 252
rect 436 248 456 249
rect 440 244 456 248
rect 436 243 456 244
rect 419 229 471 230
rect 423 225 435 229
rect 439 225 451 229
rect 455 225 471 229
rect 419 224 471 225
rect 431 217 435 224
rect 457 221 461 224
rect 423 180 426 197
rect 448 183 452 186
rect 423 178 442 180
rect 322 160 374 164
rect 423 177 431 178
rect 435 177 442 178
rect 290 154 294 160
rect 290 150 310 154
rect 377 49 381 174
rect 423 170 427 174
rect 391 166 423 170
rect 431 170 435 174
rect 439 163 442 177
rect 449 164 452 183
rect 482 186 486 269
rect 459 174 512 178
rect 455 170 459 174
rect 439 161 444 163
rect 423 158 444 161
rect 449 160 459 164
rect 423 147 426 158
rect 449 157 452 160
rect 448 152 452 157
rect 431 130 435 137
rect 457 130 461 137
rect 419 129 471 130
rect 423 125 435 129
rect 439 125 451 129
rect 455 125 471 129
rect 419 124 471 125
rect 508 49 512 174
rect 517 -18 521 367
rect 387 -22 521 -18
rect 387 -34 391 -22
<< m2contact >>
rect 336 416 340 420
rect 328 406 332 410
rect 370 426 374 430
rect 435 426 439 430
rect 121 174 125 178
rect 175 174 179 178
rect 131 166 135 170
rect 203 160 207 164
rect 408 412 412 416
rect 377 406 381 410
rect 453 412 457 416
rect 478 367 482 371
rect 517 367 521 371
rect 444 269 448 273
rect 482 269 486 273
rect 290 160 294 164
rect 377 174 381 178
rect 431 174 435 178
rect 387 166 391 170
rect 482 182 486 186
rect 459 160 463 164
<< metal2 >>
rect 374 426 435 430
rect 312 416 336 420
rect 412 412 453 416
rect 332 406 377 410
rect 482 367 517 371
rect 448 269 482 273
rect 125 174 175 178
rect 381 174 431 178
rect 131 -18 135 166
rect 207 160 290 164
rect 387 48 391 166
rect 482 164 486 182
rect 463 160 486 164
rect 387 -18 391 45
rect 131 -22 391 -18
rect 255 -35 259 -22
<< m1p >>
rect 427 422 431 426
rect 435 422 439 426
rect 459 422 463 426
rect 336 412 340 416
rect 459 412 463 416
rect 328 402 332 406
rect 448 279 452 283
rect 440 269 444 273
rect 423 170 427 174
rect 431 170 435 174
rect 455 170 459 174
rect 455 160 459 164
use MUX2X1  MUX2X1_0
timestamp 1053021328
transform 1 0 165 0 1 127
box -5 -3 53 105
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 308 0 1 127
box -9 -3 26 105
use shift_lut_slice  shift_lut_slice_0
array 0 3 128 0 0 108
timestamp 1382949514
transform 1 0 8 0 1 0
box -8 0 120 108
<< labels >>
rlabel metal1 425 172 425 172 1 S
rlabel metal1 425 227 425 227 6 vdd
rlabel metal1 425 127 425 127 8 gnd
rlabel metal1 457 162 457 162 1 Y
rlabel metal1 457 172 457 172 1 A
rlabel metal1 433 172 433 172 1 B
rlabel metal1 442 271 442 271 6 A
rlabel metal1 450 281 450 281 6 Y
rlabel metal1 442 346 442 346 6 vdd
rlabel metal1 442 246 442 246 8 gnd
rlabel metal1 429 424 429 424 1 S
rlabel metal1 429 479 429 479 6 vdd
rlabel metal1 429 379 429 379 8 gnd
rlabel metal1 461 414 461 414 1 Y
rlabel metal1 461 424 461 424 1 A
rlabel metal1 437 424 437 424 1 B
rlabel metal1 387 -34 391 -30 0 B
rlabel metal2 255 -35 259 -31 0 A
rlabel metal2 312 416 316 420 0 F
rlabel metal1 330 379 330 379 8 gnd
rlabel metal1 330 479 330 479 6 vdd
rlabel metal1 338 414 338 414 6 Y
rlabel metal1 330 404 330 404 6 A
<< end >>
