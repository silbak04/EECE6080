magic
tech scmos
timestamp 1383633248
<< error_s >>
rect 1170 49 1172 52
rect 1757 49 1759 52
rect 1173 46 1175 49
rect 1760 46 1762 49
<< error_ps >>
rect 583 162 585 165
rect 586 159 588 162
rect 583 49 585 52
rect 586 46 588 49
<< m2contact >>
rect 919 -69 923 -65
rect 1019 -70 1023 -66
rect 1119 -70 1123 -66
rect 1219 -70 1223 -66
rect 1319 -70 1323 -66
rect 1419 -70 1423 -66
rect 1519 -70 1523 -66
rect 1619 -70 1623 -66
<< metal2 >>
rect 528 228 1173 232
rect 449 217 453 226
rect 1169 219 1173 228
rect 449 214 582 217
rect 1116 116 2347 119
rect 450 105 453 113
rect 525 112 529 115
rect 525 109 595 112
rect 450 102 582 105
rect 592 104 595 109
rect 1036 110 1040 113
rect 1152 110 1760 112
rect 1036 109 1760 110
rect 1036 107 1155 109
rect 1169 104 1173 106
rect 1756 105 1760 109
rect 2343 106 2347 116
rect 592 103 1173 104
rect 592 102 1170 103
rect 592 101 1169 102
rect 449 -22 453 5
rect 525 -10 529 5
rect 1036 -1 1040 0
rect 1112 -1 1116 0
rect 1036 -4 1106 -1
rect 1112 -4 1223 -1
rect 1623 -3 1627 0
rect 1102 -9 1106 -4
rect 525 -13 1023 -10
rect 1102 -13 1123 -9
rect 449 -25 923 -22
rect 919 -65 923 -25
rect 1019 -66 1023 -13
rect 1119 -66 1123 -13
rect 1219 -66 1223 -4
rect 1319 -6 1627 -3
rect 1319 -66 1323 -6
rect 1699 -9 1703 0
rect 1419 -12 1703 -9
rect 1419 -66 1422 -12
rect 2210 -19 2214 0
rect 1519 -23 2214 -19
rect 1519 -66 1522 -23
rect 2287 -29 2290 0
rect 1619 -33 2290 -29
rect 1619 -66 1623 -33
use lut  lut_2
timestamp 1383530834
transform 1 0 -2 0 1 226
box 0 0 593 108
use lut  lut_1
array 0 1 587 0 0 108
timestamp 1383530834
transform 1 0 -2 0 1 113
box 0 0 593 108
use lut  lut_0
array 0 3 587 0 0 108
timestamp 1383530834
transform 1 0 -2 0 1 0
box 0 0 593 108
use p_shifter  p_shifter_0
timestamp 1383633248
transform 1 0 821 0 1 -113
box -36 0 812 108
<< end >>
