magic
tech scmos
timestamp 1384162313
<< metal1 >>
rect 1498 684 1524 687
rect 2335 614 2339 620
rect 2336 501 2339 507
rect 508 341 511 375
rect 515 347 518 409
rect 1739 388 1749 394
rect 2335 388 2339 394
rect 1739 362 1745 388
rect 1132 356 1745 362
rect 515 344 1148 347
rect 508 338 1142 341
rect 1139 267 1142 338
rect 1145 274 1148 344
rect 1145 271 2383 274
rect 1139 264 2389 267
rect 1105 257 2395 260
rect 1099 250 2401 253
<< m2contact >>
rect 1524 692 1528 696
rect 1524 684 1528 688
rect 2335 536 2339 540
rect 2335 423 2339 427
rect 514 409 518 413
rect 508 375 512 379
rect 2335 310 2339 314
rect 2383 271 2387 275
rect 2389 264 2393 268
rect 1101 257 1105 261
rect 2395 257 2399 261
rect 1095 250 1099 254
rect 2401 250 2405 254
<< metal2 >>
rect 1528 693 2429 696
rect 1528 684 2423 687
rect 2339 571 2417 574
rect 2339 536 2411 540
rect 1167 517 1172 519
rect -82 495 1165 498
rect -82 489 1159 492
rect -82 483 1153 486
rect -82 477 1147 480
rect -82 471 1141 474
rect -82 465 1135 468
rect -82 456 1126 459
rect -82 450 545 453
rect -82 444 538 447
rect 502 432 524 435
rect 511 409 514 412
rect 521 353 524 432
rect 535 405 538 444
rect 542 440 545 450
rect 1132 439 1135 465
rect 1120 436 1135 439
rect 1138 409 1141 471
rect 1120 406 1141 409
rect 535 402 542 405
rect 1144 379 1147 477
rect 1150 385 1153 483
rect 1156 427 1159 489
rect 1162 457 1165 495
rect 2339 458 2405 461
rect 1156 424 1163 427
rect 2339 423 2399 427
rect 1150 382 1752 385
rect 1144 376 1746 379
rect 990 353 994 357
rect 1070 356 1154 359
rect 521 350 994 353
rect 1094 296 1104 300
rect 1095 254 1098 266
rect 1101 261 1104 296
rect 1150 292 1154 356
rect 1743 314 1746 376
rect 1749 344 1752 382
rect 2339 345 2393 348
rect 1743 311 1749 314
rect 2339 310 2387 314
rect 1150 288 1754 292
rect 2384 275 2387 310
rect 2390 268 2393 345
rect 2396 261 2399 423
rect 2402 254 2405 458
rect 2408 186 2411 536
rect 2272 183 2411 186
rect 2269 155 2272 156
rect 2414 155 2417 571
rect 2269 152 2417 155
rect 2420 73 2423 684
rect 2210 70 2423 73
rect 2426 12 2429 693
rect 1532 9 2429 12
use lut  lut_0
timestamp 1384162313
transform 1 0 539 0 1 356
box 0 0 593 108
use tree  tree_1
timestamp 1384162313
transform -1 0 2340 0 -1 620
box -2 -113 2352 334
use tree  tree_0
timestamp 1384162313
transform 1 0 -80 0 1 103
box -2 -113 2352 334
<< end >>
