magic
tech scmos
timestamp 1384231894
<< metal1 >>
rect 37 36 51 40
rect 47 26 51 36
use MUX2X1  MUX2X1_0
timestamp 1384231894
transform 1 0 3 0 1 3
box -5 -5 53 105
use INVX1  INVX1_0
timestamp 1384231894
transform 1 0 45 0 1 3
box -9 -5 26 105
<< end >>
