magic
tech scmos
timestamp 1384152407
<< metal1 >>
rect 325 2038 338 2050
rect -1006 2029 -708 2038
rect -699 2029 792 2038
rect 801 2029 1092 2038
rect 1101 2029 1692 2038
rect 1701 2029 1968 2038
rect -1006 -928 -997 2029
rect -977 2012 -462 2020
rect -986 2011 -462 2012
rect -453 2011 -408 2020
rect -399 2011 -108 2020
rect -99 2011 492 2020
rect 501 2011 1038 2020
rect 1047 2011 1338 2020
rect 1347 2011 1392 2020
rect 1401 2011 1940 2020
rect -986 1578 -978 2011
rect 1633 1697 1931 1703
rect -969 1672 -741 1678
rect -145 1673 -142 1694
rect -123 1676 -75 1679
rect -739 1622 -736 1662
rect 1526 1642 1534 1645
rect 1632 1643 1645 1647
rect -124 1622 -93 1625
rect 1940 1603 1948 2011
rect 1634 1597 1948 1603
rect -986 1572 -736 1578
rect -986 1309 -978 1572
rect -127 1566 -114 1569
rect -986 1303 87 1309
rect -986 1196 -978 1303
rect 883 1203 1930 1209
rect 1940 1196 1948 1597
rect 1959 1439 1968 2029
rect -986 1190 -642 1196
rect 1709 1193 1948 1196
rect 1709 1190 1940 1193
rect -986 911 -978 1190
rect -969 1090 -642 1096
rect 1711 1090 1931 1096
rect 1940 1083 1948 1184
rect 1959 1139 1968 1430
rect 1709 1077 1948 1083
rect -119 1032 -90 1038
rect -969 1005 -711 1011
rect -119 1005 -113 1032
rect 1711 977 1931 983
rect 1940 970 1948 1077
rect 1709 964 1948 970
rect -122 945 -119 951
rect -986 905 -706 911
rect -986 870 -978 905
rect -969 892 -711 898
rect 1940 893 1948 964
rect 1711 864 1931 870
rect -986 798 -978 861
rect 469 826 475 829
rect -850 805 -846 819
rect -986 792 -706 798
rect -986 685 -978 792
rect -969 779 -711 785
rect 1642 779 1931 785
rect 1940 685 1948 884
rect 1959 839 1968 1130
rect -986 679 -706 685
rect 1642 679 1948 685
rect -986 570 -978 679
rect -709 625 -706 672
rect -600 671 -594 679
rect 917 666 1931 672
rect -700 612 -694 638
rect -969 606 -541 612
rect 74 603 106 606
rect -761 586 -542 590
rect -986 512 -978 561
rect -761 552 -525 555
rect 67 513 70 575
rect 74 532 77 603
rect 1940 593 1948 679
rect 1940 572 1948 584
rect 917 566 1948 572
rect 1940 550 1948 566
rect 1952 560 1956 613
rect 883 544 1948 550
rect -986 506 -536 512
rect 67 510 87 513
rect -986 270 -978 506
rect 87 504 90 507
rect -755 499 -701 502
rect -97 499 -80 502
rect -850 482 -846 494
rect -837 482 -833 494
rect -755 490 -701 493
rect 883 444 1931 450
rect 1940 437 1948 544
rect 1959 539 1968 830
rect 1971 580 1975 1386
rect 1709 431 1948 437
rect 1711 331 1931 337
rect 1940 324 1948 431
rect 1709 318 1948 324
rect 1940 293 1948 318
rect -986 152 -978 261
rect -125 273 -90 279
rect -125 252 -119 273
rect -969 246 -742 252
rect 1711 218 1931 224
rect 1940 211 1948 284
rect 1959 239 1968 530
rect 1709 205 1948 211
rect -745 192 -738 196
rect -122 186 -119 192
rect -986 146 -742 152
rect -986 39 -978 146
rect -969 133 -740 139
rect 1711 105 1931 111
rect -745 79 -738 82
rect 469 67 475 70
rect -986 33 -742 39
rect -986 -30 -978 33
rect -969 20 -741 26
rect 1642 20 1931 26
rect 1940 -7 1948 205
rect -747 -33 -737 -30
rect -986 -74 -978 -39
rect 1940 -74 1948 -16
rect -986 -80 -740 -74
rect 1642 -80 1948 -74
rect -986 -84 -978 -80
rect -986 -90 -741 -84
rect -986 -330 -978 -90
rect 917 -93 1931 -87
rect -747 -123 -738 -120
rect -816 -133 -807 -130
rect 73 -147 86 -143
rect -833 -156 -821 -152
rect -969 -179 -756 -173
rect -763 -184 -756 -179
rect -975 -190 -966 -186
rect -975 -201 -971 -190
rect -850 -220 -846 -189
rect -816 -189 -807 -186
rect -830 -214 -827 -189
rect -763 -190 -740 -184
rect -816 -197 -807 -194
rect -816 -205 -807 -202
rect 60 -214 63 -205
rect -830 -217 63 -214
rect 73 -220 77 -147
rect 117 -148 132 -145
rect 1940 -187 1948 -80
rect 917 -193 1948 -187
rect -850 -224 77 -220
rect -986 -607 -978 -339
rect -968 -513 -752 -507
rect -732 -513 -536 -507
rect -548 -567 -522 -564
rect -441 -567 -429 -563
rect -736 -577 -724 -574
rect -540 -577 -528 -573
rect -474 -576 -456 -573
rect -763 -587 -748 -583
rect -748 -601 -747 -597
rect -986 -613 -752 -607
rect -733 -613 -537 -607
rect -986 -909 -978 -613
rect 1940 -909 1948 -193
rect -986 -917 -983 -909
rect -972 -917 -708 -909
rect -697 -917 -408 -909
rect -399 -917 -108 -909
rect -99 -917 438 -909
rect 446 -917 1038 -909
rect 1047 -917 1092 -909
rect 1101 -917 1338 -909
rect 1347 -917 1392 -909
rect 1401 -917 1638 -909
rect 1647 -917 1692 -909
rect 1701 -917 1938 -909
rect 1947 -917 1948 -909
rect 628 -921 640 -917
rect 1959 -928 1968 230
rect 1972 215 1975 543
rect -1006 -937 -462 -928
rect -453 -937 192 -928
rect 201 -937 792 -928
rect 801 -937 1968 -928
rect 628 -950 640 -945
rect 628 -956 635 -950
<< m2contact >>
rect -708 2029 -699 2038
rect 792 2029 801 2038
rect 1092 2029 1101 2038
rect 1692 2029 1701 2038
rect -986 2012 -977 2020
rect -462 2011 -453 2020
rect -408 2011 -399 2020
rect -108 2011 -99 2020
rect 492 2011 501 2020
rect 1038 2011 1047 2020
rect 1338 2011 1347 2020
rect 1392 2011 1401 2020
rect 1940 2011 1948 2020
rect -997 1672 -991 1678
rect -145 1694 -141 1698
rect 1931 1697 1937 1703
rect -975 1672 -969 1678
rect -127 1676 -123 1680
rect -75 1676 -71 1680
rect -145 1669 -141 1673
rect -739 1662 -735 1666
rect 1522 1642 1526 1646
rect 1645 1643 1649 1647
rect -128 1622 -124 1626
rect -93 1622 -89 1626
rect 1953 1697 1959 1703
rect -131 1565 -127 1569
rect -114 1565 -110 1569
rect 1930 1203 1936 1209
rect 1959 1430 1968 1439
rect 1953 1203 1959 1209
rect -997 1090 -991 1096
rect -997 1005 -991 1011
rect 1940 1184 1948 1193
rect -975 1090 -969 1096
rect 1931 1090 1937 1096
rect 1959 1130 1968 1139
rect 1953 1090 1959 1096
rect -975 1005 -969 1011
rect 1931 977 1937 983
rect 1953 977 1959 983
rect -997 892 -991 898
rect -975 892 -969 898
rect 1940 884 1948 893
rect -986 861 -978 870
rect 1931 864 1937 870
rect -850 819 -846 823
rect -850 801 -846 805
rect -997 779 -991 785
rect -975 779 -969 785
rect 1931 779 1937 785
rect 1953 864 1959 870
rect 1959 830 1968 839
rect 1953 779 1959 785
rect -997 606 -991 612
rect -709 672 -705 676
rect 1931 666 1937 672
rect -634 655 -630 659
rect -644 639 -640 643
rect -709 621 -705 625
rect -975 606 -969 612
rect 128 611 132 615
rect -765 586 -761 590
rect -542 586 -538 590
rect -986 561 -978 570
rect 67 575 71 579
rect -765 552 -761 556
rect 1953 666 1959 672
rect 1940 584 1948 593
rect 1952 613 1956 617
rect 1952 556 1956 560
rect 74 528 78 532
rect -759 499 -755 503
rect -701 499 -697 503
rect -101 498 -97 502
rect -80 498 -76 502
rect -850 494 -846 498
rect -850 478 -846 482
rect -837 494 -833 498
rect -759 490 -755 494
rect -701 490 -697 494
rect -837 478 -833 482
rect 1931 444 1937 450
rect 1971 1386 1975 1390
rect 1971 576 1975 580
rect 1959 530 1968 539
rect 1953 444 1959 450
rect 1931 331 1937 337
rect 1953 331 1959 337
rect 1940 284 1948 293
rect -986 261 -978 270
rect -997 246 -991 252
rect -975 246 -969 252
rect 1931 218 1937 224
rect 1972 543 1976 547
rect 1959 230 1969 239
rect 1953 218 1959 224
rect -749 192 -745 196
rect -722 182 -718 186
rect -997 133 -991 139
rect -975 133 -969 139
rect 1931 105 1937 111
rect -749 79 -745 83
rect -722 69 -718 73
rect -997 20 -991 26
rect -975 20 -969 26
rect 1931 20 1937 26
rect 1953 105 1959 111
rect 1953 20 1959 26
rect 1940 -16 1948 -7
rect -986 -39 -978 -30
rect -751 -34 -747 -30
rect -722 -44 -718 -40
rect -997 -179 -991 -173
rect 1931 -93 1937 -87
rect -751 -123 -747 -119
rect -630 -120 -626 -116
rect -820 -134 -816 -130
rect -807 -134 -803 -130
rect -720 -134 -716 -130
rect -696 -134 -692 -130
rect -688 -134 -684 -130
rect -680 -134 -676 -130
rect -672 -134 -668 -130
rect -648 -134 -644 -130
rect -837 -156 -833 -152
rect -821 -156 -817 -152
rect -975 -179 -969 -173
rect -966 -190 -962 -186
rect -850 -189 -846 -185
rect -975 -205 -971 -201
rect -830 -189 -826 -185
rect -820 -189 -816 -185
rect -807 -189 -803 -185
rect -820 -197 -816 -193
rect -807 -197 -803 -193
rect -820 -205 -816 -201
rect -807 -205 -803 -201
rect 60 -205 64 -201
rect 113 -148 117 -144
rect 1953 -93 1959 -87
rect -986 -339 -978 -330
rect -997 -513 -991 -507
rect -974 -513 -968 -507
rect -552 -567 -548 -563
rect -429 -567 -425 -563
rect -724 -577 -720 -573
rect -544 -577 -540 -573
rect -456 -576 -452 -572
rect -767 -587 -763 -583
rect -983 -919 -972 -909
rect -708 -918 -697 -909
rect -408 -917 -399 -909
rect -108 -917 -99 -909
rect 438 -917 446 -909
rect 1038 -917 1047 -909
rect 1092 -917 1101 -909
rect 1338 -917 1347 -909
rect 1392 -917 1401 -909
rect 1638 -917 1647 -909
rect 1692 -917 1701 -909
rect 1938 -917 1947 -909
rect 628 -925 640 -921
rect 1972 211 1976 215
rect -462 -937 -453 -928
rect 192 -937 201 -928
rect 792 -937 801 -928
rect 628 -945 640 -941
<< metal2 >>
rect -1008 2044 -999 2050
rect -975 2044 -966 2053
rect -1008 2041 -966 2044
rect -986 2020 -977 2041
rect -762 2010 -753 2050
rect -708 2038 -699 2051
rect -762 2005 -746 2010
rect -991 1672 -975 1678
rect -751 1656 -746 2005
rect -675 2008 -666 2050
rect -462 2020 -453 2050
rect -408 2020 -399 2052
rect -375 2020 -366 2051
rect -399 2011 -366 2020
rect -162 2018 -153 2050
rect -108 2020 -99 2051
rect -75 2020 -66 2050
rect -162 2011 -133 2018
rect -99 2011 -66 2020
rect -675 2004 -142 2008
rect -145 1698 -142 2004
rect -138 2000 -133 2011
rect 138 2006 147 2050
rect 492 2020 501 2050
rect 525 2020 534 2050
rect 501 2011 534 2020
rect 738 2007 747 2050
rect 792 2038 801 2050
rect 825 2009 834 2050
rect 1038 2020 1047 2050
rect 1092 2038 1101 2052
rect -136 1685 -133 2000
rect -739 1682 -133 1685
rect -120 2003 147 2006
rect 167 2003 747 2007
rect 753 2006 834 2009
rect 1125 2010 1134 2050
rect 1338 2020 1347 2051
rect 1392 2020 1401 2051
rect 1425 2020 1434 2051
rect 1401 2011 1434 2020
rect -739 1666 -736 1682
rect -158 1676 -127 1679
rect -145 1656 -142 1669
rect -751 1652 -733 1656
rect -623 1652 -614 1656
rect -151 1652 -142 1656
rect -152 1622 -128 1625
rect -291 1561 -287 1572
rect -215 1569 -211 1578
rect -215 1566 -131 1569
rect -120 1561 -117 2003
rect 167 1841 173 2003
rect -100 1838 173 1841
rect -100 1569 -97 1838
rect 753 1831 756 2006
rect 1125 1848 1135 2010
rect 1638 2008 1647 2050
rect 1692 2038 1701 2051
rect 1725 2009 1734 2051
rect 1938 2020 1947 2050
rect -81 1828 756 1831
rect 771 1846 1135 1848
rect 1522 2005 1647 2008
rect 1689 2005 1734 2009
rect 771 1845 1133 1846
rect -81 1625 -78 1828
rect 771 1824 774 1845
rect -74 1821 774 1824
rect -74 1680 -71 1821
rect 1522 1646 1525 2005
rect 1689 1844 1692 2005
rect 1670 1840 1692 1844
rect 1670 1647 1674 1840
rect 1937 1697 1953 1703
rect 1649 1643 1674 1647
rect -89 1622 -78 1625
rect -110 1566 -97 1569
rect -291 1558 -117 1561
rect 1968 1430 1981 1439
rect 1971 1397 1988 1406
rect 1971 1390 1975 1397
rect 739 1309 824 1312
rect 63 1302 1806 1306
rect 63 1290 66 1302
rect -819 1287 79 1290
rect -1019 1111 -969 1116
rect -1019 1107 -846 1111
rect -991 1090 -975 1096
rect -991 1005 -975 1011
rect -1019 894 -1006 903
rect -1010 870 -1006 894
rect -991 892 -975 898
rect -1019 861 -986 870
rect -850 823 -846 1107
rect -1021 813 -978 816
rect -1021 808 -833 813
rect -1021 807 -978 808
rect -991 779 -975 785
rect -991 606 -975 612
rect -1020 594 -978 602
rect -986 570 -978 594
rect -1019 561 -986 570
rect -1019 507 -992 516
rect -996 491 -992 507
rect -850 498 -846 801
rect -837 498 -833 808
rect -996 487 -850 491
rect -846 487 -826 491
rect -1019 294 -978 303
rect -986 270 -978 294
rect -1019 261 -986 270
rect -991 246 -975 252
rect -1019 207 -963 216
rect -991 133 -975 139
rect -991 20 -975 26
rect -1019 -6 -978 3
rect -986 -30 -978 -6
rect -1019 -39 -986 -30
rect -1019 -93 -1011 -84
rect -1014 -193 -1011 -93
rect -991 -179 -975 -173
rect -966 -186 -963 207
rect -850 -185 -846 478
rect -837 -152 -833 478
rect -830 -185 -826 487
rect -819 -130 -816 1287
rect -813 1263 87 1266
rect -820 -185 -817 -156
rect -1014 -197 -820 -193
rect -971 -205 -820 -201
rect -813 -208 -810 1263
rect -807 1122 -641 1125
rect -807 66 -804 1122
rect -801 1112 -640 1115
rect -801 82 -798 1112
rect 1803 1104 1806 1302
rect 1936 1203 1953 1209
rect 1948 1184 1981 1193
rect 1968 1130 1982 1139
rect 1969 1104 1986 1106
rect 1803 1101 1986 1104
rect 1969 1097 1986 1101
rect 1937 1090 1953 1096
rect -795 1071 -711 1074
rect -795 179 -792 1071
rect -789 1065 -712 1068
rect -789 195 -786 1065
rect -783 1059 -712 1062
rect -783 264 -780 1059
rect -777 1053 -704 1056
rect -777 270 -774 1053
rect -771 1047 -711 1050
rect -771 555 -768 1047
rect -765 1041 -710 1044
rect -765 590 -762 1041
rect -758 1032 -711 1035
rect 532 1033 535 1039
rect -771 552 -765 555
rect -758 503 -755 1032
rect -752 1026 -712 1029
rect -758 276 -755 490
rect -752 285 -749 1026
rect -746 1020 -710 1023
rect -699 1020 -696 1023
rect -746 291 -743 1020
rect -740 985 -708 988
rect -740 297 -737 985
rect 502 982 508 985
rect 1937 977 1953 983
rect -734 951 -708 954
rect -734 303 -731 951
rect 1119 920 1122 926
rect 1948 884 1981 893
rect -728 872 -708 875
rect -728 309 -725 872
rect 1937 864 1953 870
rect -722 838 -709 841
rect -722 315 -719 838
rect 1968 830 1981 839
rect 1972 797 1983 806
rect 1937 779 1953 785
rect -716 760 -708 763
rect -716 659 -712 760
rect 1642 728 1647 731
rect -709 676 -706 725
rect 1937 666 1953 672
rect -716 655 -634 659
rect 66 654 75 657
rect 923 646 932 650
rect -644 634 -640 639
rect -716 630 -640 634
rect -716 357 -713 630
rect -709 390 -706 621
rect 1972 617 1975 797
rect 46 609 63 612
rect 1956 613 1975 617
rect 50 586 57 590
rect 54 560 57 586
rect 60 569 63 609
rect 129 579 132 611
rect 1948 584 1982 593
rect 71 576 132 579
rect 1778 576 1971 580
rect 1778 569 1781 576
rect 60 566 1781 569
rect 54 556 1952 560
rect 48 550 51 556
rect 48 547 1781 550
rect 1778 539 1781 547
rect 1953 543 1972 546
rect 1953 539 1956 543
rect 1778 536 1956 539
rect 1968 530 1982 539
rect -697 499 -101 502
rect -91 493 -87 506
rect -15 502 -11 506
rect 1972 502 1982 506
rect -76 499 -11 502
rect 1803 499 1982 502
rect -697 490 -87 493
rect 68 466 77 470
rect -709 387 -639 390
rect -716 353 -642 357
rect -722 312 -711 315
rect -728 306 -712 309
rect -734 300 -710 303
rect -740 294 -712 297
rect -746 288 -709 291
rect -752 282 -711 285
rect -758 273 -712 276
rect 532 274 535 280
rect -777 267 -708 270
rect -783 261 -690 264
rect -722 226 -709 230
rect -789 192 -749 195
rect -722 186 -718 226
rect 502 223 508 226
rect -709 179 -706 192
rect -795 176 -706 179
rect 1119 161 1122 167
rect -722 114 -703 117
rect -722 113 -709 114
rect -801 79 -749 82
rect -722 73 -718 113
rect -709 66 -706 79
rect -807 63 -706 66
rect -722 0 -708 4
rect -751 -119 -748 -34
rect -722 -40 -719 0
rect 1642 -31 1647 -28
rect -709 -77 -706 -34
rect -709 -80 -627 -77
rect -630 -116 -627 -80
rect 923 -113 932 -109
rect -803 -133 -720 -130
rect -696 -186 -693 -134
rect -803 -189 -693 -186
rect -684 -194 -680 -130
rect -803 -197 -680 -194
rect -672 -202 -669 -134
rect -803 -205 -669 -202
rect -648 -208 -645 -134
rect 60 -142 116 -139
rect 60 -201 63 -142
rect 113 -144 116 -142
rect 1803 -207 1806 499
rect 1972 497 1982 499
rect 1937 444 1953 450
rect 1937 331 1953 337
rect 1948 284 1983 293
rect 1969 230 1981 239
rect 1937 218 1953 224
rect 1972 206 1976 211
rect 1972 197 1981 206
rect 1937 105 1953 111
rect 1937 20 1953 26
rect 1948 -16 1981 -7
rect 1937 -93 1953 -87
rect 1147 -208 1806 -207
rect -813 -211 1806 -208
rect 1147 -212 1806 -211
rect -1020 -306 -978 -297
rect -986 -330 -978 -306
rect -1019 -339 -986 -330
rect -991 -513 -974 -507
rect -425 -567 -412 -563
rect -720 -577 -580 -573
rect -767 -904 -764 -587
rect -767 -909 -753 -904
rect -584 -906 -580 -577
rect -552 -903 -548 -567
rect -452 -576 -428 -573
rect -544 -735 -540 -577
rect -432 -728 -428 -576
rect -416 -718 -412 -567
rect -416 -722 886 -718
rect -432 -731 291 -728
rect -544 -739 8 -735
rect -552 -906 -153 -903
rect -675 -909 -580 -906
rect -1008 -919 -983 -909
rect -972 -919 -966 -909
rect -1008 -951 -999 -919
rect -975 -950 -966 -919
rect -762 -951 -753 -909
rect -708 -950 -699 -918
rect -675 -950 -666 -909
rect -399 -917 -366 -910
rect -462 -951 -453 -937
rect -408 -950 -399 -917
rect -375 -951 -366 -917
rect -162 -951 -153 -906
rect -99 -917 -67 -909
rect -108 -950 -99 -917
rect -76 -951 -67 -917
rect -4 -923 8 -739
rect 288 -902 291 -731
rect 225 -907 291 -902
rect 882 -903 886 -722
rect 825 -907 886 -903
rect -4 -926 145 -923
rect 138 -950 145 -926
rect 192 -950 201 -937
rect 225 -950 234 -907
rect 438 -951 446 -917
rect 628 -941 640 -925
rect 628 -950 640 -945
rect 792 -951 800 -937
rect 825 -951 834 -907
rect 1038 -951 1047 -917
rect 1101 -917 1134 -909
rect 1092 -956 1101 -917
rect 1125 -956 1134 -917
rect 1338 -956 1347 -917
rect 1401 -917 1434 -909
rect 1392 -956 1401 -917
rect 1425 -957 1434 -917
rect 1638 -956 1647 -917
rect 1701 -917 1734 -909
rect 1692 -956 1701 -917
rect 1725 -956 1734 -917
rect 1938 -958 1947 -917
<< m1p >>
rect -128 1622 -124 1626
rect -93 1622 -89 1626
use lut  lut_1
timestamp 1383979221
transform 1 0 -742 0 1 1572
box 0 0 593 108
use shift_slice  shift_slice_0
timestamp 1383130333
transform 1 0 1527 0 1 1597
box 0 0 112 108
use BUFX4  BUFX4_4
timestamp 1053722803
transform 0 -1 -597 1 0 637
box -9 -3 37 105
use lut_p_tree  lut_p_tree_1
timestamp 1384142942
transform 1 0 -630 0 1 576
box -82 -10 2429 733
use lut  lut_0
timestamp 1383979221
transform 1 0 -542 0 1 506
box 0 0 593 108
use BUFX4  BUFX4_3
timestamp 1053722803
transform 1 0 -740 0 1 149
box -9 -3 37 105
use BUFX4  BUFX4_2
timestamp 1053722803
transform 1 0 -740 0 1 36
box -9 -3 37 105
use BUFX4  BUFX4_0
timestamp 1053722803
transform 1 0 -740 0 1 -77
box -9 -3 37 105
use mux  mux_0
timestamp 1382957000
transform -1 0 -679 0 -1 -84
box -2 0 71 108
use mux  mux_1
timestamp 1382957000
transform 1 0 -685 0 -1 -84
box -2 0 71 108
use BUFX4  BUFX4_1
timestamp 1053722803
transform 1 0 84 0 1 -190
box -9 -3 37 105
use lut_p_tree  lut_p_tree_0
timestamp 1384142942
transform 1 0 -630 0 1 -183
box -82 -10 2429 733
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 -750 0 1 -610
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_0
timestamp 1383129201
transform 1 0 -535 0 1 -610
box -8 -3 104 105
<< labels >>
rlabel m2contact -820 -205 -816 -201 0 L_IN
rlabel metal2 73 -142 77 -139 0 P_IN
rlabel metal2 1778 576 1781 580 0 F
rlabel metal1 1959 2029 1968 2038 0 VDD
rlabel metal2 79 1263 87 1266 0 P_OUT
rlabel metal2 -630 -84 -627 -80 0 M2
rlabel metal2 -751 -119 -748 -115 0 M1
rlabel m2contact 1940 2011 1948 2020 0 GND
rlabel metal2 923 -113 932 -109 0 PQ0
rlabel metal2 68 466 77 470 0 PQ1
rlabel metal2 923 646 932 650 0 PQ2
rlabel metal2 1642 -31 1647 -28 0 LO_0
rlabel metal2 1642 728 1647 731 0 LO_2
rlabel metal2 -647 1122 -642 1125 0 LO_3
rlabel metal1 469 67 475 70 0 LO_4
rlabel metal2 532 274 535 280 0 LO_5
rlabel metal1 469 826 475 829 0 LO_6
rlabel metal2 532 1033 535 1039 0 LO_7
rlabel metal1 -122 186 -119 192 0 LO_8
rlabel metal2 1119 161 1122 167 0 LO_9
rlabel metal2 1119 920 1122 926 0 LO_11
rlabel metal1 -122 945 -119 951 0 LO_10
rlabel metal2 502 223 508 226 0 LO_12
rlabel metal2 502 982 508 985 0 LO_13
rlabel metal2 1778 536 1781 540 0 L_OUT
rlabel m2contact -820 -197 -816 -193 0 TMEI
rlabel m2contact -820 -189 -816 -185 0 LCLKI
rlabel metal1 73 -147 77 -143 0 PCLKI
rlabel metal2 66 654 75 657 0 PQ2_1
rlabel metal2 -651 387 -642 390 0 LO_1
<< end >>
