magic
tech scmos
timestamp 1383038773
use DFFPOSX1  DFFPOSX1_0
array 0 15 97 0 0 108
timestamp 1383038773
transform 1 0 8 0 1 3
box -8 -3 104 105
<< end >>
