magic
tech scmos
timestamp 1380881990
<< ntransistor >>
rect -44 20 -40 22
rect 86 20 90 22
rect -44 3 -40 5
rect 86 2 90 4
rect -44 -17 -40 -15
rect 86 -16 90 -14
rect 86 -34 90 -32
rect -44 -43 -40 -41
rect 29 -54 33 -52
rect -44 -61 -40 -59
rect 86 -54 90 -52
rect 29 -74 33 -72
rect 86 -74 90 -72
rect -44 -95 -40 -93
rect 29 -94 33 -92
rect 86 -97 90 -95
rect -44 -113 -40 -111
<< ptransistor >>
rect -28 20 -24 22
rect 102 20 106 22
rect -28 3 -24 5
rect 102 2 106 4
rect -28 -17 -24 -15
rect 102 -16 106 -14
rect 102 -34 106 -32
rect -23 -43 -19 -41
rect 13 -54 17 -52
rect -23 -61 -19 -59
rect 102 -54 106 -52
rect 13 -74 17 -72
rect 102 -74 106 -72
rect -16 -95 -12 -93
rect 13 -94 17 -92
rect 102 -97 106 -95
rect -16 -113 -12 -111
<< ndiffusion >>
rect -44 22 -40 23
rect 86 22 90 24
rect -44 19 -40 20
rect 86 18 90 20
rect -44 5 -40 7
rect -44 -1 -40 3
rect 86 4 90 6
rect 86 0 90 2
rect -44 -15 -40 -13
rect 86 -14 90 -12
rect -44 -19 -40 -17
rect 86 -18 90 -16
rect -44 -41 -40 -37
rect 86 -32 90 -30
rect -44 -45 -40 -43
rect 86 -36 90 -34
rect -44 -59 -40 -57
rect 29 -52 33 -50
rect -44 -63 -40 -61
rect 29 -58 33 -54
rect 86 -52 90 -48
rect 86 -56 90 -54
rect 29 -72 33 -70
rect 86 -72 90 -68
rect 29 -76 33 -74
rect 86 -76 90 -74
rect -44 -93 -40 -89
rect -44 -97 -40 -95
rect 29 -92 33 -88
rect 29 -96 33 -94
rect 86 -95 90 -94
rect 86 -98 90 -97
rect -44 -111 -40 -109
rect -44 -117 -40 -113
<< pdiffusion >>
rect -28 22 -24 23
rect 102 22 106 24
rect -28 19 -24 20
rect 102 18 106 20
rect -28 5 -24 7
rect -28 -1 -24 3
rect 102 4 106 6
rect 102 0 106 2
rect -28 -15 -24 -13
rect 102 -14 106 -12
rect -28 -19 -24 -17
rect 102 -18 106 -16
rect 102 -32 106 -30
rect -23 -41 -19 -35
rect 102 -36 106 -34
rect -23 -45 -19 -43
rect 13 -52 17 -50
rect -23 -59 -19 -57
rect 13 -58 17 -54
rect -23 -63 -19 -61
rect 102 -52 106 -48
rect 102 -56 106 -54
rect 13 -72 17 -70
rect 102 -72 106 -68
rect 13 -76 17 -74
rect 102 -76 106 -74
rect -16 -93 -12 -89
rect 13 -92 17 -88
rect -16 -97 -12 -95
rect 13 -96 17 -94
rect 102 -95 106 -94
rect 102 -98 106 -97
rect -16 -111 -12 -109
rect -16 -117 -12 -113
<< ndcontact >>
rect -44 23 -40 27
rect 86 24 90 28
rect -44 15 -40 19
rect 86 14 90 18
rect -44 7 -40 11
rect 86 6 90 10
rect -44 -5 -40 -1
rect 86 -4 90 0
rect -44 -13 -40 -9
rect 86 -12 90 -8
rect -44 -23 -40 -19
rect 86 -22 90 -18
rect 86 -30 90 -26
rect -44 -37 -40 -33
rect 86 -40 90 -36
rect -44 -49 -40 -45
rect -44 -57 -40 -53
rect 29 -50 33 -46
rect 86 -48 90 -44
rect -44 -67 -40 -63
rect 29 -62 33 -58
rect 86 -60 90 -56
rect 29 -70 33 -66
rect 86 -68 90 -64
rect 29 -80 33 -76
rect 86 -80 90 -76
rect -44 -89 -40 -85
rect 29 -88 33 -84
rect 86 -94 90 -90
rect -44 -101 -40 -97
rect 29 -100 33 -96
rect 86 -102 90 -98
rect -44 -109 -40 -105
rect -44 -121 -40 -117
<< pdcontact >>
rect -28 23 -24 27
rect 102 24 106 28
rect -28 15 -24 19
rect 102 14 106 18
rect -28 7 -24 11
rect 102 6 106 10
rect -28 -5 -24 -1
rect 102 -4 106 0
rect -28 -13 -24 -9
rect 102 -12 106 -8
rect -28 -23 -24 -19
rect 102 -22 106 -18
rect -23 -35 -19 -31
rect 102 -30 106 -26
rect 102 -40 106 -36
rect -23 -49 -19 -45
rect 13 -50 17 -46
rect -23 -57 -19 -53
rect 13 -62 17 -58
rect 102 -48 106 -44
rect 102 -60 106 -56
rect -23 -67 -19 -63
rect 13 -70 17 -66
rect 102 -68 106 -64
rect 13 -80 17 -76
rect 102 -80 106 -76
rect -16 -89 -12 -85
rect 13 -88 17 -84
rect -16 -101 -12 -97
rect 13 -100 17 -96
rect 102 -94 106 -90
rect 102 -102 106 -98
rect -16 -109 -12 -105
rect -16 -121 -12 -117
<< polysilicon >>
rect -46 20 -44 22
rect -40 20 -28 22
rect -24 20 86 22
rect 90 20 102 22
rect 106 20 124 22
rect -68 3 -44 5
rect -40 3 -36 5
rect -32 3 -28 5
rect -24 3 -22 5
rect 48 2 86 4
rect 90 2 102 4
rect 106 2 108 4
rect -47 -17 -44 -15
rect -40 -17 -28 -15
rect -24 -17 -22 -15
rect 84 -16 86 -14
rect 90 -16 102 -14
rect 106 -16 108 -14
rect 62 -34 86 -32
rect 90 -34 102 -32
rect 106 -34 108 -32
rect -47 -43 -44 -41
rect -40 -43 -37 -41
rect -33 -43 -23 -41
rect -19 -43 65 -41
rect 69 -43 124 -41
rect -4 -54 13 -52
rect 17 -54 29 -52
rect 33 -54 35 -52
rect -54 -61 -44 -59
rect -40 -61 -23 -59
rect -19 -61 -17 -59
rect 83 -54 86 -52
rect 90 -54 102 -52
rect 106 -54 108 -52
rect -4 -74 13 -72
rect 17 -74 29 -72
rect 33 -74 35 -72
rect 84 -74 86 -72
rect 90 -74 102 -72
rect 106 -74 109 -72
rect -47 -95 -44 -93
rect -40 -95 -37 -93
rect -33 -95 -16 -93
rect -12 -95 -10 -93
rect 10 -94 13 -92
rect 17 -94 29 -92
rect 33 -94 35 -92
rect 83 -97 86 -95
rect 90 -97 102 -95
rect 106 -97 108 -95
rect -68 -113 -44 -111
rect -40 -113 -34 -111
rect -30 -113 -16 -111
rect -12 -113 -10 -111
<< polycontact >>
rect -72 2 -68 6
rect -36 2 -32 6
rect 44 1 48 5
rect -51 -18 -47 -14
rect 94 -14 98 -10
rect 58 -35 62 -31
rect -37 -44 -33 -40
rect 65 -44 69 -40
rect -58 -62 -54 -58
rect -8 -55 -4 -51
rect 79 -55 83 -51
rect -8 -75 -4 -71
rect 109 -75 113 -71
rect -51 -96 -47 -92
rect -37 -96 -33 -92
rect 6 -95 10 -91
rect 79 -98 83 -94
rect -72 -114 -68 -110
rect -34 -114 -30 -110
<< metal1 >>
rect -65 27 -61 31
rect -1 27 3 31
rect -65 23 -44 27
rect -24 23 3 27
rect -65 11 -61 23
rect -40 15 -28 19
rect -65 7 -44 11
rect -72 -110 -68 2
rect -65 -33 -61 7
rect -36 6 -32 15
rect -1 11 3 23
rect -24 7 3 11
rect -44 -9 -40 -5
rect -36 -5 -28 -1
rect -51 -26 -47 -18
rect -36 -19 -32 -5
rect -1 -9 3 7
rect -24 -13 3 -9
rect -40 -23 -28 -19
rect -24 -23 -20 -19
rect -51 -30 -33 -26
rect -65 -37 -44 -33
rect -65 -85 -61 -37
rect -37 -40 -33 -30
rect -30 -38 -26 -23
rect -1 -26 3 -13
rect -23 -30 3 -26
rect -23 -31 -19 -30
rect -30 -42 -4 -38
rect -44 -53 -40 -49
rect -30 -49 -23 -45
rect -58 -78 -54 -62
rect -30 -63 -26 -49
rect -8 -51 -4 -42
rect -19 -57 -11 -53
rect -1 -46 3 -30
rect 29 -33 33 35
rect 21 -37 33 -33
rect -1 -50 13 -46
rect -14 -58 -11 -57
rect -1 -58 3 -50
rect 21 -58 25 -37
rect 37 -46 41 35
rect 33 -50 41 -46
rect 44 5 48 35
rect -14 -62 3 -58
rect 17 -62 25 -58
rect -40 -67 -23 -63
rect -23 -71 -19 -67
rect -1 -66 3 -62
rect -1 -70 13 -66
rect -23 -75 -8 -71
rect -58 -82 -33 -78
rect -16 -79 -12 -75
rect -65 -89 -44 -85
rect -65 -128 -61 -89
rect -37 -92 -33 -82
rect -1 -84 3 -70
rect 21 -76 25 -62
rect 29 -66 33 -62
rect 17 -80 25 -76
rect -1 -85 13 -84
rect -12 -88 13 -85
rect -12 -89 3 -88
rect -51 -124 -47 -96
rect -44 -105 -40 -101
rect -23 -101 -16 -97
rect -23 -117 -19 -101
rect -1 -105 3 -89
rect -12 -109 3 -105
rect 6 -117 10 -95
rect 21 -96 25 -80
rect 29 -84 33 -80
rect 44 -94 48 1
rect 51 16 55 35
rect 116 28 120 32
rect 72 24 86 28
rect 106 24 120 28
rect 72 16 76 24
rect 51 12 76 16
rect 51 -86 55 12
rect 72 -8 76 12
rect 86 10 90 14
rect 94 14 102 18
rect 94 0 98 14
rect 116 10 120 24
rect 106 6 120 10
rect 90 -4 102 0
rect 72 -12 86 -8
rect 94 -10 98 -4
rect 116 -8 120 6
rect 58 -76 62 -35
rect 65 -51 69 -44
rect 72 -44 76 -12
rect 106 -12 120 -8
rect 86 -26 90 -22
rect 79 -36 83 -26
rect 94 -22 102 -18
rect 94 -36 98 -22
rect 116 -26 120 -12
rect 106 -30 120 -26
rect 79 -40 86 -36
rect 90 -40 102 -36
rect 116 -44 120 -30
rect 72 -48 86 -44
rect 106 -48 120 -44
rect 65 -55 79 -51
rect 86 -64 90 -60
rect 94 -60 102 -56
rect 94 -76 98 -60
rect 116 -64 120 -48
rect 106 -68 120 -64
rect 58 -80 86 -76
rect 90 -80 102 -76
rect 109 -83 113 -75
rect 51 -90 90 -86
rect 94 -87 113 -83
rect 17 -100 29 -96
rect 44 -98 79 -94
rect 94 -98 98 -87
rect 116 -90 120 -68
rect 106 -94 120 -90
rect -40 -121 -16 -117
rect -12 -121 10 -117
rect 13 -107 33 -103
rect 13 -124 17 -107
rect -51 -128 17 -124
rect 29 -128 33 -107
rect 44 -128 48 -98
rect 90 -102 102 -98
rect 116 -128 120 -94
<< labels >>
rlabel metal1 79 -30 83 -26 0 MUX_OUT
rlabel polysilicon 120 20 124 22 0 A
rlabel polysilicon 120 -43 124 -41 0 B
rlabel metal1 44 -128 48 -124 0 SEL
rlabel metal1 51 31 55 35 0 GND
rlabel metal1 44 31 48 35 0 SEL
rlabel metal1 37 31 41 35 0 GND
rlabel metal1 29 -128 33 -124 0 C_IN
rlabel metal1 29 31 33 35 0 C_OUT
rlabel metal1 -24 -23 -20 -19 0 A_OUT
rlabel metal1 -16 -79 -12 -75 0 B_OUT
rlabel metal1 -4 -121 0 -117 0 CIN_OUT
rlabel metal1 -1 27 3 31 0 VDD
rlabel metal1 -65 27 -61 31 0 GND
rlabel metal1 116 28 120 32 0 VDD
<< end >>
