magic
tech scmos
timestamp 1383556561
<< metal1 >>
rect -755 1020 -739 1023
rect 87 612 115 615
rect -761 587 -525 590
rect -761 552 -525 555
rect 87 507 90 612
rect 94 603 108 606
rect 94 532 97 603
rect 87 503 104 507
rect -755 499 -701 502
rect -82 499 -65 502
rect -755 490 -701 493
<< m2contact >>
rect -759 1019 -755 1023
rect -739 1019 -735 1023
rect -765 587 -761 591
rect -525 586 -521 590
rect -765 552 -761 556
rect 94 528 98 532
rect -759 499 -755 503
rect -701 499 -697 503
rect -86 498 -82 502
rect -65 498 -61 502
rect -759 490 -755 494
rect -701 490 -697 494
<< metal2 >>
rect -807 1122 -641 1125
rect -807 83 -804 1122
rect -801 1112 -640 1115
rect -801 117 -798 1112
rect -795 1071 -711 1074
rect -795 195 -792 1071
rect -789 1065 -712 1068
rect -789 230 -786 1065
rect -783 1059 -712 1062
rect -783 264 -780 1059
rect -777 1053 -704 1056
rect -777 270 -774 1053
rect -771 1047 -711 1050
rect -771 555 -768 1047
rect -765 1041 -710 1044
rect -765 591 -762 1041
rect -752 1032 -711 1035
rect -771 552 -765 555
rect -758 503 -755 1019
rect -758 276 -755 490
rect -752 285 -749 1032
rect -746 1026 -712 1029
rect -746 291 -743 1026
rect -735 1020 -696 1023
rect -740 985 -708 988
rect -740 297 -737 985
rect -734 951 -708 954
rect -734 303 -731 951
rect -728 872 -708 875
rect -728 309 -725 872
rect -722 838 -709 841
rect -722 315 -719 838
rect -716 760 -708 763
rect -716 357 -713 760
rect -709 388 -706 725
rect 61 609 81 612
rect 66 587 74 590
rect 71 559 74 587
rect 78 569 81 609
rect 78 566 1761 569
rect 71 556 1761 559
rect 63 550 66 556
rect 63 547 1761 550
rect -697 499 -86 502
rect -76 493 -72 506
rect 0 502 4 507
rect -61 499 4 502
rect -697 490 -72 493
rect -709 385 -639 388
rect -716 354 -642 357
rect -722 312 -711 315
rect -728 306 -712 309
rect -734 300 -710 303
rect -740 294 -712 297
rect -746 288 -709 291
rect -752 282 -711 285
rect -758 273 -712 276
rect -777 267 -708 270
rect -783 261 -690 264
rect -789 227 -708 230
rect -795 192 -709 195
rect -801 114 -703 117
rect -807 80 -709 83
use lut_p_tree  lut_p_tree_1
timestamp 1383549043
transform 1 0 -630 0 1 576
box -82 -10 2393 733
use lut  lut_0
timestamp 1383530834
transform 1 0 -527 0 1 506
box 0 0 593 108
use lut_p_tree  lut_p_tree_0
timestamp 1383549043
transform 1 0 -630 0 1 -183
box -82 -10 2393 733
<< end >>
