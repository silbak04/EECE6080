magic
tech scmos
timestamp 1382962255
use box  box_0
timestamp 1382962255
transform 1 0 1396 0 1 1153
box -166 109 2354 2621
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1072203966
transform 1 0 -4 0 1 0
box 4 0 5004 5000
<< end >>
