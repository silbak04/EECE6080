* SPICE3 file created from part_5b.ext - technology: scmos

.option scale=0.3u

M1000 GND A0 part_5_0[0]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=1856 pd=1504 as=20 ps=18 
M1001 VDD A0 part_5_0[0]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=3584 pd=2880 as=20 ps=18 
M1002 GND A0 part_5_0[0]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1003 VDD A0 part_5_0[0]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1004 GND part_5_0[0]/a_n72_n114# part_5_0[0]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1005 VDD part_5_0[0]/a_n72_n114# part_5_0[0]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1006 part_5_0[0]/a_86_4# part_5_0[0]/SEL part_5_0[0]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1007 VDD part_5_0[0]/SEL part_5_0[0]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1008 part_5_0[0]/a_n44_n15# B0 part_5_0[0]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1009 VDD B0 part_5_0[0]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1010 GND part_5_0[0]/a_84_n16# part_5_0[0]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1011 VDD part_5_0[0]/a_84_n16# F0 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1012 part_5_0[0]/a_86_n32# part_5_0[0]/a_58_n35# F0 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1013 VDD part_5_0[0]/a_58_n35# F0 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1014 GND B0 part_5_0[0]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1015 VDD B0 part_5_0[0]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1016 VDD part_5_0[0]/A_OUT part_5_0[1]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1017 GND part_5_0[0]/A_OUT part_5_0[0]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1018 part_5_0[0]/a_n44_n59# GND part_5_0[0]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1019 VDD GND part_5_0[0]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1020 GND B0 part_5_0[0]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1021 VDD B0 part_5_0[0]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1022 VDD part_5_0[0]/B_OUT part_5_0[1]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1023 part_5_0[0]/a_29_n72# part_5_0[0]/B_OUT part_5_0[0]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1024 part_5_0[0]/a_86_n72# part_5_0[0]/a_84_n74# part_5_0[0]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1025 VDD part_5_0[0]/a_84_n74# part_5_0[0]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1026 GND GND part_5_0[0]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1027 VDD GND part_5_0[0]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1028 VDD part_5_0[0]/CIN_OUT part_5_0[1]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1029 part_5_0[0]/a_29_n92# part_5_0[0]/CIN_OUT part_5_0[1]/C_IN Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1030 GND part_5_0[0]/SEL part_5_0[0]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1031 VDD part_5_0[0]/SEL part_5_0[0]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1032 part_5_0[0]/a_n44_n111# part_5_0[0]/a_n72_n114# part_5_0[0]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1033 VDD part_5_0[0]/a_n72_n114# part_5_0[0]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1034 GND A1 part_5_0[1]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1035 VDD A1 part_5_0[1]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1036 GND A1 part_5_0[1]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1037 VDD A1 part_5_0[1]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1038 GND part_5_0[1]/a_n72_n114# part_5_0[1]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1039 VDD part_5_0[1]/a_n72_n114# part_5_0[1]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1040 part_5_0[1]/a_86_4# part_5_0[0]/SEL part_5_0[1]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1041 VDD part_5_0[0]/SEL part_5_0[1]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1042 part_5_0[1]/a_n44_n15# B1 part_5_0[1]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1043 VDD B1 part_5_0[1]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1044 GND part_5_0[1]/a_84_n16# part_5_0[1]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1045 VDD part_5_0[1]/a_84_n16# F1 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1046 part_5_0[1]/a_86_n32# part_5_0[1]/a_58_n35# F1 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1047 VDD part_5_0[1]/a_58_n35# F1 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1048 GND B1 part_5_0[1]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1049 VDD B1 part_5_0[1]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1050 VDD part_5_0[1]/A_OUT part_5_0[2]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1051 GND part_5_0[1]/A_OUT part_5_0[1]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1052 part_5_0[1]/a_n44_n59# part_5_0[1]/C_IN part_5_0[1]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1053 VDD part_5_0[1]/C_IN part_5_0[1]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1054 GND B1 part_5_0[1]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1055 VDD B1 part_5_0[1]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1056 VDD part_5_0[1]/B_OUT part_5_0[2]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1057 part_5_0[1]/a_29_n72# part_5_0[1]/B_OUT part_5_0[1]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1058 part_5_0[1]/a_86_n72# part_5_0[1]/a_84_n74# part_5_0[1]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1059 VDD part_5_0[1]/a_84_n74# part_5_0[1]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1060 GND part_5_0[1]/C_IN part_5_0[1]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1061 VDD part_5_0[1]/C_IN part_5_0[1]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1062 VDD part_5_0[1]/CIN_OUT part_5_0[2]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1063 part_5_0[1]/a_29_n92# part_5_0[1]/CIN_OUT part_5_0[2]/C_IN Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1064 GND part_5_0[0]/SEL part_5_0[1]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1065 VDD part_5_0[0]/SEL part_5_0[1]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1066 part_5_0[1]/a_n44_n111# part_5_0[1]/a_n72_n114# part_5_0[1]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1067 VDD part_5_0[1]/a_n72_n114# part_5_0[1]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1068 GND A2 part_5_0[2]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1069 VDD A2 part_5_0[2]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1070 GND A2 part_5_0[2]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1071 VDD A2 part_5_0[2]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1072 GND part_5_0[2]/a_n72_n114# part_5_0[2]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1073 VDD part_5_0[2]/a_n72_n114# part_5_0[2]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1074 part_5_0[2]/a_86_4# part_5_0[0]/SEL part_5_0[2]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1075 VDD part_5_0[0]/SEL part_5_0[2]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1076 part_5_0[2]/a_n44_n15# B2 part_5_0[2]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1077 VDD B2 part_5_0[2]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1078 GND part_5_0[2]/a_84_n16# part_5_0[2]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1079 VDD part_5_0[2]/a_84_n16# F2 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1080 part_5_0[2]/a_86_n32# part_5_0[2]/a_58_n35# F2 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1081 VDD part_5_0[2]/a_58_n35# F2 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1082 GND B2 part_5_0[2]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1083 VDD B2 part_5_0[2]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1084 VDD part_5_0[2]/A_OUT part_5_0[3]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1085 GND part_5_0[2]/A_OUT part_5_0[2]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1086 part_5_0[2]/a_n44_n59# part_5_0[2]/C_IN part_5_0[2]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1087 VDD part_5_0[2]/C_IN part_5_0[2]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1088 GND B2 part_5_0[2]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1089 VDD B2 part_5_0[2]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1090 VDD part_5_0[2]/B_OUT part_5_0[3]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1091 part_5_0[2]/a_29_n72# part_5_0[2]/B_OUT part_5_0[2]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1092 part_5_0[2]/a_86_n72# part_5_0[2]/a_84_n74# part_5_0[2]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1093 VDD part_5_0[2]/a_84_n74# part_5_0[2]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1094 GND part_5_0[2]/C_IN part_5_0[2]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1095 VDD part_5_0[2]/C_IN part_5_0[2]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1096 VDD part_5_0[2]/CIN_OUT part_5_0[3]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1097 part_5_0[2]/a_29_n92# part_5_0[2]/CIN_OUT part_5_0[3]/C_IN Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1098 GND part_5_0[0]/SEL part_5_0[2]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1099 VDD part_5_0[0]/SEL part_5_0[2]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1100 part_5_0[2]/a_n44_n111# part_5_0[2]/a_n72_n114# part_5_0[2]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1101 VDD part_5_0[2]/a_n72_n114# part_5_0[2]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1102 GND A3 part_5_0[3]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1103 VDD A3 part_5_0[3]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1104 GND A3 part_5_0[3]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1105 VDD A3 part_5_0[3]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1106 GND part_5_0[3]/a_n72_n114# part_5_0[3]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1107 VDD part_5_0[3]/a_n72_n114# part_5_0[3]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1108 part_5_0[3]/a_86_4# part_5_0[0]/SEL part_5_0[3]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1109 VDD part_5_0[0]/SEL part_5_0[3]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1110 part_5_0[3]/a_n44_n15# B3 part_5_0[3]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1111 VDD B3 part_5_0[3]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1112 GND part_5_0[3]/a_84_n16# part_5_0[3]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1113 VDD part_5_0[3]/a_84_n16# F3 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1114 part_5_0[3]/a_86_n32# part_5_0[3]/a_58_n35# F3 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1115 VDD part_5_0[3]/a_58_n35# F3 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1116 GND B3 part_5_0[3]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1117 VDD B3 part_5_0[3]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1118 VDD part_5_0[3]/A_OUT part_5_0[4]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1119 GND part_5_0[3]/A_OUT part_5_0[3]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1120 part_5_0[3]/a_n44_n59# part_5_0[3]/C_IN part_5_0[3]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1121 VDD part_5_0[3]/C_IN part_5_0[3]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1122 GND B3 part_5_0[3]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1123 VDD B3 part_5_0[3]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1124 VDD part_5_0[3]/B_OUT part_5_0[4]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1125 part_5_0[3]/a_29_n72# part_5_0[3]/B_OUT part_5_0[3]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1126 part_5_0[3]/a_86_n72# part_5_0[3]/a_84_n74# part_5_0[3]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1127 VDD part_5_0[3]/a_84_n74# part_5_0[3]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1128 GND part_5_0[3]/C_IN part_5_0[3]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1129 VDD part_5_0[3]/C_IN part_5_0[3]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1130 VDD part_5_0[3]/CIN_OUT part_5_0[4]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1131 part_5_0[3]/a_29_n92# part_5_0[3]/CIN_OUT part_5_0[4]/C_IN Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1132 GND part_5_0[0]/SEL part_5_0[3]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1133 VDD part_5_0[0]/SEL part_5_0[3]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1134 part_5_0[3]/a_n44_n111# part_5_0[3]/a_n72_n114# part_5_0[3]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1135 VDD part_5_0[3]/a_n72_n114# part_5_0[3]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1136 GND A4 part_5_0[4]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1137 VDD A4 part_5_0[4]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1138 GND A4 part_5_0[4]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1139 VDD A4 part_5_0[4]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1140 GND part_5_0[4]/a_n72_n114# part_5_0[4]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1141 VDD part_5_0[4]/a_n72_n114# part_5_0[4]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1142 part_5_0[4]/a_86_4# part_5_0[0]/SEL part_5_0[4]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1143 VDD part_5_0[0]/SEL part_5_0[4]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1144 part_5_0[4]/a_n44_n15# B4 part_5_0[4]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1145 VDD B4 part_5_0[4]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1146 GND part_5_0[4]/a_84_n16# part_5_0[4]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1147 VDD part_5_0[4]/a_84_n16# F4 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1148 part_5_0[4]/a_86_n32# part_5_0[4]/a_58_n35# F4 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1149 VDD part_5_0[4]/a_58_n35# F4 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1150 GND B4 part_5_0[4]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1151 VDD B4 part_5_0[4]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1152 VDD part_5_0[4]/A_OUT part_5_0[5]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1153 GND part_5_0[4]/A_OUT part_5_0[4]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1154 part_5_0[4]/a_n44_n59# part_5_0[4]/C_IN part_5_0[4]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1155 VDD part_5_0[4]/C_IN part_5_0[4]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1156 GND B4 part_5_0[4]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1157 VDD B4 part_5_0[4]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1158 VDD part_5_0[4]/B_OUT part_5_0[5]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1159 part_5_0[4]/a_29_n72# part_5_0[4]/B_OUT part_5_0[4]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1160 part_5_0[4]/a_86_n72# part_5_0[4]/a_84_n74# part_5_0[4]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1161 VDD part_5_0[4]/a_84_n74# part_5_0[4]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1162 GND part_5_0[4]/C_IN part_5_0[4]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1163 VDD part_5_0[4]/C_IN part_5_0[4]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1164 VDD part_5_0[4]/CIN_OUT part_5_0[5]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1165 part_5_0[4]/a_29_n92# part_5_0[4]/CIN_OUT part_5_0[5]/C_IN Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1166 GND part_5_0[0]/SEL part_5_0[4]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1167 VDD part_5_0[0]/SEL part_5_0[4]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1168 part_5_0[4]/a_n44_n111# part_5_0[4]/a_n72_n114# part_5_0[4]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1169 VDD part_5_0[4]/a_n72_n114# part_5_0[4]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1170 GND A5 part_5_0[5]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1171 VDD A5 part_5_0[5]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1172 GND A5 part_5_0[5]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1173 VDD A5 part_5_0[5]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1174 GND part_5_0[5]/a_n72_n114# part_5_0[5]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1175 VDD part_5_0[5]/a_n72_n114# part_5_0[5]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1176 part_5_0[5]/a_86_4# part_5_0[0]/SEL part_5_0[5]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1177 VDD part_5_0[0]/SEL part_5_0[5]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1178 part_5_0[5]/a_n44_n15# B5 part_5_0[5]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1179 VDD B5 part_5_0[5]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1180 GND part_5_0[5]/a_84_n16# part_5_0[5]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1181 VDD part_5_0[5]/a_84_n16# F5 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1182 part_5_0[5]/a_86_n32# part_5_0[5]/a_58_n35# F5 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1183 VDD part_5_0[5]/a_58_n35# F5 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1184 GND B5 part_5_0[5]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1185 VDD B5 part_5_0[5]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1186 VDD part_5_0[5]/A_OUT part_5_0[6]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1187 GND part_5_0[5]/A_OUT part_5_0[5]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1188 part_5_0[5]/a_n44_n59# part_5_0[5]/C_IN part_5_0[5]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1189 VDD part_5_0[5]/C_IN part_5_0[5]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1190 GND B5 part_5_0[5]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1191 VDD B5 part_5_0[5]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1192 VDD part_5_0[5]/B_OUT part_5_0[6]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1193 part_5_0[5]/a_29_n72# part_5_0[5]/B_OUT part_5_0[5]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1194 part_5_0[5]/a_86_n72# part_5_0[5]/a_84_n74# part_5_0[5]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1195 VDD part_5_0[5]/a_84_n74# part_5_0[5]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1196 GND part_5_0[5]/C_IN part_5_0[5]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1197 VDD part_5_0[5]/C_IN part_5_0[5]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1198 VDD part_5_0[5]/CIN_OUT part_5_0[6]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1199 part_5_0[5]/a_29_n92# part_5_0[5]/CIN_OUT part_5_0[6]/C_IN Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1200 GND part_5_0[0]/SEL part_5_0[5]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1201 VDD part_5_0[0]/SEL part_5_0[5]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1202 part_5_0[5]/a_n44_n111# part_5_0[5]/a_n72_n114# part_5_0[5]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1203 VDD part_5_0[5]/a_n72_n114# part_5_0[5]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1204 GND A6 part_5_0[6]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1205 VDD A6 part_5_0[6]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1206 GND A6 part_5_0[6]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1207 VDD A6 part_5_0[6]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1208 GND part_5_0[6]/a_n72_n114# part_5_0[6]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1209 VDD part_5_0[6]/a_n72_n114# part_5_0[6]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1210 part_5_0[6]/a_86_4# part_5_0[0]/SEL part_5_0[6]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1211 VDD part_5_0[0]/SEL part_5_0[6]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1212 part_5_0[6]/a_n44_n15# B6 part_5_0[6]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1213 VDD B6 part_5_0[6]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1214 GND part_5_0[6]/a_84_n16# part_5_0[6]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1215 VDD part_5_0[6]/a_84_n16# F6 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1216 part_5_0[6]/a_86_n32# part_5_0[6]/a_58_n35# F6 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1217 VDD part_5_0[6]/a_58_n35# F6 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1218 GND B6 part_5_0[6]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1219 VDD B6 part_5_0[6]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1220 VDD part_5_0[6]/A_OUT part_5_0[7]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1221 GND part_5_0[6]/A_OUT part_5_0[6]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1222 part_5_0[6]/a_n44_n59# part_5_0[6]/C_IN part_5_0[6]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1223 VDD part_5_0[6]/C_IN part_5_0[6]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1224 GND B6 part_5_0[6]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1225 VDD B6 part_5_0[6]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1226 VDD part_5_0[6]/B_OUT part_5_0[7]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1227 part_5_0[6]/a_29_n72# part_5_0[6]/B_OUT part_5_0[6]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1228 part_5_0[6]/a_86_n72# part_5_0[6]/a_84_n74# part_5_0[6]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1229 VDD part_5_0[6]/a_84_n74# part_5_0[6]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1230 GND part_5_0[6]/C_IN part_5_0[6]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1231 VDD part_5_0[6]/C_IN part_5_0[6]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1232 VDD part_5_0[6]/CIN_OUT part_5_0[7]/C_IN Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1233 part_5_0[6]/a_29_n92# part_5_0[6]/CIN_OUT part_5_0[7]/C_IN Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1234 GND part_5_0[0]/SEL part_5_0[6]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1235 VDD part_5_0[0]/SEL part_5_0[6]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1236 part_5_0[6]/a_n44_n111# part_5_0[6]/a_n72_n114# part_5_0[6]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1237 VDD part_5_0[6]/a_n72_n114# part_5_0[6]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1238 GND A7 part_5_0[7]/a_n72_n114# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1239 VDD A7 part_5_0[7]/a_n72_n114# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1240 GND A7 part_5_0[7]/a_86_4# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1241 VDD A7 part_5_0[7]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1242 GND part_5_0[7]/a_n72_n114# part_5_0[7]/a_n44_n15# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1243 VDD part_5_0[7]/a_n72_n114# part_5_0[7]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1244 part_5_0[7]/a_86_4# part_5_0[0]/SEL part_5_0[7]/a_84_n16# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1245 VDD part_5_0[0]/SEL part_5_0[7]/a_84_n16# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1246 part_5_0[7]/a_n44_n15# B7 part_5_0[7]/A_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1247 VDD B7 part_5_0[7]/A_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1248 GND part_5_0[7]/a_84_n16# part_5_0[7]/a_86_n32# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1249 VDD part_5_0[7]/a_84_n16# F7 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1250 part_5_0[7]/a_86_n32# part_5_0[7]/a_58_n35# F7 Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1251 VDD part_5_0[7]/a_58_n35# F7 Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1252 GND B7 part_5_0[7]/a_n44_n59# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1253 VDD B7 part_5_0[7]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1254 VDD part_5_0[7]/A_OUT part_5_0[0]/SEL Vdd pfet w=4 l=2
+ ad=0 pd=0 as=80 ps=64 
M1255 GND part_5_0[7]/A_OUT part_5_0[7]/a_29_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1256 part_5_0[7]/a_n44_n59# part_5_0[7]/C_IN part_5_0[7]/B_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1257 VDD part_5_0[7]/C_IN part_5_0[7]/B_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1258 GND B7 part_5_0[7]/a_86_n72# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1259 VDD B7 part_5_0[7]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1260 VDD part_5_0[7]/B_OUT part_5_0[0]/SEL Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1261 part_5_0[7]/a_29_n72# part_5_0[7]/B_OUT part_5_0[7]/a_29_n92# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1262 part_5_0[7]/a_86_n72# part_5_0[7]/a_84_n74# part_5_0[7]/a_58_n35# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1263 VDD part_5_0[7]/a_84_n74# part_5_0[7]/a_58_n35# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1264 GND part_5_0[7]/C_IN part_5_0[7]/a_n44_n111# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=48 ps=40 
M1265 VDD part_5_0[7]/C_IN part_5_0[7]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=56 ps=44 
M1266 VDD part_5_0[7]/CIN_OUT part_5_0[0]/SEL Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
M1267 part_5_0[7]/a_29_n92# part_5_0[7]/CIN_OUT part_5_0[0]/SEL Gnd nfet w=4 l=2
+ ad=0 pd=0 as=24 ps=20 
M1268 GND part_5_0[0]/SEL part_5_0[7]/a_84_n74# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1269 VDD part_5_0[0]/SEL part_5_0[7]/a_84_n74# Vdd pfet w=4 l=2
+ ad=0 pd=0 as=20 ps=18 
M1270 part_5_0[7]/a_n44_n111# part_5_0[7]/a_n72_n114# part_5_0[7]/CIN_OUT Gnd nfet w=4 l=2
+ ad=0 pd=0 as=32 ps=24 
M1271 VDD part_5_0[7]/a_n72_n114# part_5_0[7]/CIN_OUT Vdd pfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0 
C0 part_5_0[7]/CIN_OUT gnd! 5.6fF
C1 part_5_0[7]/a_84_n74# gnd! 3.3fF
C2 part_5_0[7]/C_IN gnd! 19.9fF
C3 part_5_0[7]/B_OUT gnd! 4.2fF
C4 part_5_0[7]/a_58_n35# gnd! 7.4fF
C5 part_5_0[0]/SEL gnd! 107.8fF
C6 part_5_0[7]/A_OUT gnd! 6.2fF
C7 part_5_0[7]/a_84_n16# gnd! 2.9fF
C8 part_5_0[7]/a_n72_n114# gnd! 10.2fF
C9 part_5_0[6]/CIN_OUT gnd! 5.6fF
C10 part_5_0[6]/a_84_n74# gnd! 3.3fF
C11 part_5_0[6]/C_IN gnd! 19.9fF
C12 part_5_0[6]/B_OUT gnd! 4.2fF
C13 part_5_0[6]/a_58_n35# gnd! 7.4fF
C14 part_5_0[6]/A_OUT gnd! 6.2fF
C15 part_5_0[6]/a_84_n16# gnd! 2.9fF
C16 part_5_0[6]/a_n72_n114# gnd! 10.2fF
C17 part_5_0[5]/CIN_OUT gnd! 5.6fF
C18 part_5_0[5]/a_84_n74# gnd! 3.3fF
C19 part_5_0[5]/C_IN gnd! 19.9fF
C20 part_5_0[5]/B_OUT gnd! 4.2fF
C21 part_5_0[5]/a_58_n35# gnd! 7.4fF
C22 part_5_0[5]/A_OUT gnd! 6.2fF
C23 part_5_0[5]/a_84_n16# gnd! 2.9fF
C24 part_5_0[5]/a_n72_n114# gnd! 10.2fF
C25 part_5_0[4]/CIN_OUT gnd! 5.6fF
C26 part_5_0[4]/a_84_n74# gnd! 3.3fF
C27 part_5_0[4]/C_IN gnd! 19.9fF
C28 part_5_0[4]/B_OUT gnd! 4.2fF
C29 part_5_0[4]/a_58_n35# gnd! 7.4fF
C30 part_5_0[4]/A_OUT gnd! 6.2fF
C31 part_5_0[4]/a_84_n16# gnd! 2.9fF
C32 part_5_0[4]/a_n72_n114# gnd! 10.2fF
C33 part_5_0[3]/CIN_OUT gnd! 5.6fF
C34 part_5_0[3]/a_84_n74# gnd! 3.3fF
C35 part_5_0[3]/C_IN gnd! 19.9fF
C36 part_5_0[3]/B_OUT gnd! 4.2fF
C37 part_5_0[3]/a_58_n35# gnd! 7.4fF
C38 part_5_0[3]/A_OUT gnd! 6.2fF
C39 part_5_0[3]/a_84_n16# gnd! 2.9fF
C40 part_5_0[3]/a_n72_n114# gnd! 10.2fF
C41 part_5_0[2]/CIN_OUT gnd! 5.6fF
C42 part_5_0[2]/a_84_n74# gnd! 3.3fF
C43 part_5_0[2]/C_IN gnd! 19.9fF
C44 part_5_0[2]/B_OUT gnd! 4.2fF
C45 part_5_0[2]/a_58_n35# gnd! 7.4fF
C46 part_5_0[2]/A_OUT gnd! 6.2fF
C47 part_5_0[2]/a_84_n16# gnd! 2.9fF
C48 part_5_0[2]/a_n72_n114# gnd! 10.2fF
C49 part_5_0[1]/CIN_OUT gnd! 5.6fF
C50 part_5_0[1]/a_84_n74# gnd! 3.3fF
C51 part_5_0[1]/C_IN gnd! 19.9fF
C52 part_5_0[1]/B_OUT gnd! 4.2fF
C53 part_5_0[1]/a_58_n35# gnd! 7.4fF
C54 part_5_0[1]/A_OUT gnd! 6.2fF
C55 part_5_0[1]/a_84_n16# gnd! 2.9fF
C56 part_5_0[1]/a_n72_n114# gnd! 10.2fF
C57 part_5_0[0]/CIN_OUT gnd! 5.6fF
C58 part_5_0[0]/a_84_n74# gnd! 3.3fF
C59 part_5_0[0]/B_OUT gnd! 4.4fF
C60 part_5_0[0]/a_58_n35# gnd! 7.4fF
C61 part_5_0[0]/A_OUT gnd! 6.2fF
C62 part_5_0[0]/a_84_n16# gnd! 2.9fF
C63 part_5_0[0]/a_n72_n114# gnd! 10.4fF
C64 VDD gnd! 240.3fF
