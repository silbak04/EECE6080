magic
tech scmos
timestamp 1383723055
<< error_s >>
rect 1364 1890 1365 1892
rect -638 1002 -635 1006
<< metal1 >>
rect 31 1893 35 1928
rect 882 1927 883 1929
rect 879 1904 883 1927
rect 879 1900 1225 1904
rect 1221 1897 1225 1900
rect 31 1890 486 1893
rect 31 1889 490 1890
rect -358 1876 118 1880
rect 114 1776 118 1876
rect 1727 1834 1731 1927
rect 1567 1831 1731 1834
rect 1567 1829 1570 1831
rect 104 1772 118 1776
rect 910 1826 1570 1829
rect 145 934 148 1410
rect 910 1401 913 1826
rect -118 931 148 934
rect 933 1034 946 1038
rect -343 924 -124 927
rect -343 914 -340 924
rect -233 903 -230 917
rect -224 905 -221 917
rect -127 907 -124 924
rect -118 921 -114 931
rect 274 924 601 928
rect 933 921 938 1034
rect -97 917 625 921
rect 933 918 1095 921
rect 933 917 1383 918
rect -97 891 -94 917
rect 509 910 613 913
rect -67 903 135 907
rect -67 893 -63 903
rect -224 879 -221 885
rect 142 878 145 910
rect 622 904 625 917
rect 1030 914 1383 917
rect 992 910 994 914
rect 605 886 628 890
rect 624 879 628 886
rect 990 879 994 910
<< m2contact >>
rect 27 1944 31 1948
rect 875 1944 879 1948
rect 1723 1944 1727 1948
rect 486 1890 490 1894
rect 1221 1892 1225 1897
rect -362 1876 -358 1880
rect 84 1782 88 1786
rect 144 1410 148 1414
rect 910 1397 914 1401
rect -233 917 -229 921
rect -224 917 -220 921
rect -343 910 -339 914
rect 270 924 274 928
rect 601 924 605 928
rect 962 1024 966 1028
rect -118 917 -114 921
rect -233 899 -229 903
rect -224 901 -220 905
rect -127 903 -123 907
rect 142 910 146 914
rect 505 910 509 914
rect 135 903 139 907
rect -224 885 -220 889
rect -97 887 -93 891
rect -67 889 -63 893
rect 613 909 617 913
rect 1383 914 1387 918
rect 988 910 992 914
rect 622 900 626 904
rect 601 886 605 890
rect -220 858 -216 862
rect 146 858 150 862
rect 628 858 632 862
rect 994 859 998 863
<< metal2 >>
rect -3 1948 1 1953
rect 35 1951 46 1954
rect -3 1944 27 1948
rect -362 1880 -358 1921
rect -331 1877 -328 1894
rect 43 1887 46 1951
rect 845 1948 849 1953
rect 883 1951 892 1954
rect 889 1948 892 1951
rect 1693 1948 1697 1953
rect 1731 1951 1740 1954
rect 845 1944 875 1948
rect 1693 1944 1723 1948
rect 889 1904 892 1943
rect 889 1901 1244 1904
rect 517 1887 520 1895
rect 43 1884 520 1887
rect 1241 1895 1244 1901
rect 1334 1895 1338 1896
rect 1241 1892 1338 1895
rect 1364 1895 1366 1916
rect 1221 1889 1225 1892
rect 1364 1890 1368 1895
rect 1365 1889 1368 1890
rect 1221 1885 1368 1889
rect -331 1874 -20 1877
rect -23 1861 -20 1874
rect -23 1858 80 1861
rect 77 1776 80 1858
rect 1737 1835 1740 1951
rect 1597 1834 1740 1835
rect 907 1832 1740 1834
rect 907 1831 1601 1832
rect 84 1742 88 1782
rect 78 1738 88 1742
rect 907 1427 911 1831
rect 138 1410 144 1413
rect 136 935 140 1383
rect 962 1068 972 1072
rect 962 1028 966 1068
rect -233 931 140 935
rect 535 931 714 935
rect -233 921 -230 931
rect -220 918 -118 921
rect -313 912 142 914
rect -310 910 142 912
rect 270 907 274 924
rect 535 913 539 931
rect -123 903 113 906
rect 139 903 274 907
rect -233 855 -230 899
rect -224 889 -221 901
rect 110 885 113 903
rect 601 890 605 924
rect 711 914 714 931
rect 969 926 972 1037
rect 969 922 1011 926
rect 1008 917 1011 922
rect 1008 914 1356 917
rect 617 909 695 912
rect 711 910 988 914
rect 1353 911 1356 914
rect 613 908 695 909
rect 691 904 695 908
rect 691 901 984 904
rect 622 891 625 900
rect 616 887 625 891
rect 110 882 136 885
rect -216 858 -186 862
rect -233 852 -224 855
rect -190 853 -186 858
rect 133 855 136 882
rect 150 858 180 861
rect 133 852 142 855
rect 176 853 179 858
rect 616 855 619 887
rect 632 858 662 862
rect 616 852 624 855
rect 658 853 662 858
rect 981 856 984 901
rect 998 859 1027 862
rect 1006 858 1027 859
rect 981 853 993 856
rect 1024 853 1027 858
<< m1p >>
rect 910 1397 914 1401
use top_bott_tree  top_bott_tree_1
timestamp 1383721316
transform -1 0 1016 0 -1 2799
box -775 129 1777 907
use lut  lut_6
timestamp 1383712281
transform 1 0 244 0 1 1712
box -34 0 593 108
use lut  lut_5
timestamp 1383712281
transform 1 0 241 0 1 1581
box -34 0 593 108
use lut  lut_4
timestamp 1383712281
transform 1 0 242 0 1 1454
box -34 0 593 108
use lut  lut_3
timestamp 1383712281
transform 1 0 242 0 1 1335
box -34 0 593 108
use lut  lut_2
timestamp 1383712281
transform 1 0 242 0 1 1217
box -34 0 593 108
use lut  lut_1
timestamp 1383712281
transform 1 0 240 0 1 1100
box -34 0 593 108
use new_tree  new_tree_0
timestamp 1383721316
transform 0 1 -516 -1 0 1828
box -8 -123 848 655
use lut  lut_0
timestamp 1383712281
transform 1 0 240 0 1 979
box -34 0 593 108
use new_tree  new_tree_1
timestamp 1383721316
transform 0 -1 1566 1 0 982
box -8 -123 848 655
use mux  mux_0
timestamp 1382957000
transform 1 0 -768 0 1 897
box -2 0 71 108
use mux  mux_1
timestamp 1382957000
transform 1 0 -709 0 1 897
box -2 0 71 108
use top_bott_tree  top_bott_tree_0
timestamp 1383721316
transform 1 0 9 0 1 7
box -775 129 1777 907
<< end >>
