magic
tech scmos
timestamp 1384231894
<< error_s >>
rect 3 8 4 10
rect 404 8 405 10
<< nwell >>
rect 400 51 404 108
<< pwell >>
rect 93 -2 99 3
rect 189 -2 195 3
rect 285 -2 291 3
<< metal1 >>
rect 1 100 6 106
rect 394 100 407 106
rect 585 100 593 106
rect 7 46 25 49
rect 102 46 121 49
rect 198 46 217 49
rect 294 46 313 49
rect 454 39 457 44
rect 584 40 587 93
rect 581 36 587 40
rect 394 0 407 6
rect 585 0 593 6
<< m2contact >>
rect 584 93 588 97
rect 3 46 7 50
rect 98 46 102 50
rect 194 46 198 50
rect 290 46 294 50
rect 386 46 390 50
rect 18 36 22 40
rect 114 36 118 40
rect 210 36 214 40
rect 306 36 310 40
<< metal2 >>
rect 584 97 588 106
rect 3 80 593 84
rect 18 40 22 80
rect 98 4 102 46
rect 114 40 118 80
rect 194 10 198 46
rect 210 40 214 80
rect 290 16 294 46
rect 306 40 310 80
rect 386 71 411 74
rect 505 71 593 74
rect 386 50 390 71
rect 393 65 411 68
rect 393 16 396 65
rect 290 13 396 16
rect 399 59 411 62
rect 399 10 402 59
rect 194 7 402 10
rect 405 53 411 56
rect 405 4 408 53
rect 590 50 593 71
rect 465 38 468 42
rect 98 1 408 4
rect 451 0 455 6
rect 527 0 531 6
use DFFPOSX1  DFFPOSX1_0(0)
timestamp 1384231894
transform 1 0 8 0 1 3
box -8 -5 104 105
use DFFPOSX1  DFFPOSX1_0(1)
timestamp 1384231894
transform 1 0 104 0 1 3
box -8 -5 104 105
use DFFPOSX1  DFFPOSX1_0(2)
timestamp 1384231894
transform 1 0 200 0 1 3
box -8 -5 104 105
use DFFPOSX1  DFFPOSX1_0(3)
timestamp 1384231894
transform 1 0 296 0 1 3
box -8 -5 104 105
use mux_4_to_1  mux_4_to_1_0
timestamp 1384231894
transform 1 0 404 0 1 0
box 0 -2 189 108
<< labels >>
rlabel metal2 586 101 586 101 6 F
rlabel metal1 2 103 2 103 6 VDD
rlabel metal1 591 3 591 3 6 GND
rlabel metal2 529 3 529 3 6 B
rlabel metal2 453 3 453 3 6 A
rlabel metal2 4 82 4 82 6 LCLKI
rlabel metal2 591 51 591 51 6 L_OUT
rlabel metal1 105 47 105 47 6 L3
rlabel metal1 201 47 201 47 6 L2
rlabel metal1 455 42 455 42 6 MUX1
rlabel metal2 466 41 466 41 6 INV1
rlabel m2contact 5 48 5 48 6 L_IN
<< end >>
