magic
tech scmos
timestamp 1384226059
<< metal2 >>
rect -2183 1047 -2182 1056
use box  box_0
timestamp 1384217043
transform 1 0 -1163 0 1 -114
box -1021 -958 1988 2053
use IIT_Frame_PR  IIT_Frame_PR_0
timestamp 1072203966
transform 1 0 -3186 0 1 -2064
box 4 0 5004 5000
<< end >>
