magic
tech scmos
timestamp 1383892968
<< nwell >>
rect 6 -38 234 -35
<< metal1 >>
rect 234 649 284 652
rect 115 475 118 496
rect 172 15 173 19
rect 57 -6 60 0
rect 120 5 158 8
rect 86 1 90 2
rect 169 1 173 15
rect 86 -3 173 1
rect 176 -6 179 7
rect 57 -9 179 -6
rect 234 -9 237 649
rect 281 647 284 649
rect 281 644 479 647
rect 270 627 273 642
rect 282 636 284 639
rect 302 636 452 639
rect 281 626 284 636
rect 469 634 576 637
rect 218 -12 237 -9
rect 294 -11 297 1
rect 323 -4 327 1
rect 356 2 359 562
rect 356 -1 393 2
rect 407 -4 411 17
rect 418 -3 421 8
rect 323 -8 411 -4
rect 538 -5 541 3
rect 568 1 572 2
rect 568 -2 610 1
rect 647 -3 650 8
rect 657 5 661 15
rect 632 -5 650 -3
rect 538 -6 650 -5
rect 418 -11 421 -6
rect 538 -8 636 -6
rect 294 -14 421 -11
rect 482 -11 535 -10
rect 640 -11 661 -10
rect 482 -13 661 -11
rect 532 -14 643 -13
<< m2contact >>
rect 115 496 119 500
rect 115 471 119 475
rect 173 32 177 36
rect 56 0 60 4
rect 86 2 90 6
rect 116 5 120 9
rect 158 5 162 9
rect 176 7 180 11
rect 214 -12 218 -8
rect 270 642 274 646
rect 479 644 483 648
rect 278 636 282 640
rect 298 636 302 640
rect 452 636 456 640
rect 270 623 274 627
rect 465 634 469 638
rect 576 634 580 638
rect 281 622 285 626
rect 289 615 293 619
rect 296 599 300 603
rect 356 562 360 566
rect 293 1 297 5
rect 323 1 327 5
rect 415 31 419 35
rect 661 32 665 36
rect 393 -1 397 3
rect 418 8 422 12
rect 646 8 650 12
rect 538 3 542 7
rect 568 2 572 6
rect 606 1 610 5
rect 657 1 661 5
rect 478 -13 482 -9
rect 661 -13 665 -9
rect 134 -77 138 -73
rect 234 -77 238 -73
rect 334 -77 338 -73
rect 434 -77 438 -73
rect 534 -77 538 -73
rect 634 -77 638 -73
rect 734 -77 738 -73
rect 834 -77 838 -73
<< metal2 >>
rect 270 649 284 652
rect 270 646 273 649
rect 281 647 284 649
rect 281 644 301 647
rect 298 640 301 644
rect 173 636 278 639
rect 173 628 176 636
rect 203 630 293 633
rect 203 629 207 630
rect 229 623 270 626
rect 280 597 284 622
rect 289 619 293 630
rect 415 628 418 654
rect 445 630 449 655
rect 300 599 326 602
rect 280 594 292 597
rect 323 594 326 599
rect 115 566 123 569
rect 356 566 365 569
rect 115 500 118 566
rect 93 489 123 493
rect 331 489 366 492
rect -8 142 7 145
rect -8 -40 -5 142
rect 6 66 10 70
rect 6 -34 9 66
rect 93 22 96 489
rect 99 471 115 474
rect 99 28 102 471
rect 226 143 244 146
rect 99 25 139 28
rect 93 19 131 22
rect 112 9 120 13
rect 128 -28 131 19
rect 136 -22 139 25
rect 166 25 169 42
rect 204 36 207 42
rect 177 33 207 36
rect 166 22 179 25
rect 176 11 179 22
rect 158 -9 161 5
rect 158 -12 214 -9
rect 226 -16 229 143
rect 234 67 244 70
rect 234 -10 237 67
rect 331 57 334 489
rect 452 70 455 636
rect 479 637 482 644
rect 580 634 605 637
rect 465 625 469 634
rect 479 145 482 634
rect 602 568 605 634
rect 717 622 728 625
rect 602 565 611 568
rect 725 567 728 622
rect 725 564 735 567
rect 575 489 611 493
rect 479 142 491 145
rect 452 67 488 70
rect 330 31 334 57
rect 445 43 448 45
rect 330 -4 333 31
rect 408 26 411 43
rect 445 35 449 43
rect 419 32 449 35
rect 408 23 421 26
rect 418 12 421 23
rect 349 9 403 12
rect 330 -7 367 -4
rect 234 -13 359 -10
rect 226 -19 351 -16
rect 136 -25 344 -22
rect 128 -31 337 -28
rect 234 -34 237 -31
rect 6 -37 237 -34
rect -8 -43 137 -40
rect 134 -73 137 -43
rect 234 -73 237 -37
rect 334 -73 337 -31
rect 341 -38 344 -25
rect 348 -30 351 -19
rect 355 -22 359 -13
rect 364 -16 367 -7
rect 394 -10 397 -1
rect 400 -3 403 9
rect 400 -5 541 -3
rect 575 -5 578 489
rect 723 488 734 491
rect 647 39 657 42
rect 647 12 650 39
rect 691 36 695 41
rect 665 32 695 36
rect 594 9 603 12
rect 600 -2 603 9
rect 610 1 657 5
rect 723 -2 726 488
rect 600 -5 728 -2
rect 400 -6 578 -5
rect 534 -8 578 -6
rect 394 -13 478 -10
rect 364 -19 651 -16
rect 355 -25 637 -22
rect 348 -34 538 -30
rect 341 -41 437 -38
rect 434 -73 437 -41
rect 534 -73 537 -34
rect 634 -73 637 -25
rect 647 -34 651 -19
rect 661 -26 664 -13
rect 661 -29 837 -26
rect 647 -38 737 -34
rect 734 -73 737 -38
rect 834 -73 837 -29
<< m1p >>
rect 115 496 119 500
rect 115 471 119 475
rect 434 -77 438 -73
use lut  lut_0
timestamp 1383712281
transform 0 1 6 -1 0 597
box -34 0 593 108
use lut  lut_1
timestamp 1383712281
transform 0 1 123 1 0 38
box -34 0 593 108
use lut  lut_2
timestamp 1383712281
transform 0 1 243 -1 0 597
box -34 0 593 108
use lut  lut_3
timestamp 1383712281
transform 0 1 365 1 0 38
box -34 0 593 108
use lut  lut_4
timestamp 1383712281
transform 0 1 488 -1 0 597
box -34 0 593 108
use lut  lut_5
timestamp 1383712281
transform 0 1 611 1 0 38
box -34 0 593 108
use lut  lut_6
timestamp 1383712281
transform 0 1 734 1 0 36
box -34 0 593 108
use p_shifter  p_shifter_0
timestamp 1383647763
transform 1 0 36 0 1 -123
box -36 0 812 108
<< end >>
