magic
tech scmos
timestamp 1382962255
use tree  tree_2
timestamp 1382962255
transform -1 0 2186 0 -1 2604
box -2 0 2352 334
use tree  tree_1
timestamp 1382962255
transform 0 -1 2344 1 0 269
box -2 0 2352 334
use tree  tree_0
timestamp 1382962255
transform 1 0 2 0 1 122
box -2 0 2352 334
use tree  tree_3
timestamp 1382962255
transform 0 1 -161 -1 0 2461
box -2 0 2352 334
<< end >>
